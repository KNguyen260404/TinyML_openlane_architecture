VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Random_forest_top_ver2
  CLASS BLOCK ;
  FOREIGN Random_forest_top_ver2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 317.195 BY 327.915 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 13.720 10.640 16.720 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 43.720 10.640 46.720 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 73.720 10.640 76.720 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 103.720 10.640 106.720 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 133.720 10.640 136.720 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 163.720 10.640 166.720 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 193.720 10.640 196.720 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 223.720 10.640 226.720 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 253.720 10.640 256.720 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 283.720 10.640 286.720 315.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 19.080 311.660 22.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 49.080 311.660 52.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 79.080 311.660 82.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 109.080 311.660 112.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 139.080 311.660 142.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 169.080 311.660 172.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 199.080 311.660 202.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 229.080 311.660 232.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 259.080 311.660 262.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 289.080 311.660 292.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 9.020 10.640 12.020 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 39.020 10.640 42.020 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 69.020 10.640 72.020 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 99.020 10.640 102.020 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 129.020 10.640 132.020 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 159.020 10.640 162.020 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 189.020 10.640 192.020 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 219.020 10.640 222.020 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 249.020 10.640 252.020 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 279.020 10.640 282.020 315.760 ;
    END
    PORT
      LAYER met4 ;
        RECT 309.020 10.640 312.020 315.760 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 14.380 312.020 17.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 44.380 312.020 47.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 74.380 312.020 77.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 104.380 312.020 107.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 134.380 312.020 137.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 164.380 312.020 167.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 194.380 312.020 197.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 224.380 312.020 227.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 254.380 312.020 257.380 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 284.380 312.020 287.380 ;
    END
  END VPWR
  PIN arbitration_id[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.050 323.915 12.330 327.915 ;
    END
  END arbitration_id[0]
  PIN arbitration_id[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.050 323.915 35.330 327.915 ;
    END
  END arbitration_id[10]
  PIN arbitration_id[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 37.350 323.915 37.630 327.915 ;
    END
  END arbitration_id[11]
  PIN arbitration_id[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 39.650 323.915 39.930 327.915 ;
    END
  END arbitration_id[12]
  PIN arbitration_id[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 323.915 42.230 327.915 ;
    END
  END arbitration_id[13]
  PIN arbitration_id[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 44.250 323.915 44.530 327.915 ;
    END
  END arbitration_id[14]
  PIN arbitration_id[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 46.550 323.915 46.830 327.915 ;
    END
  END arbitration_id[15]
  PIN arbitration_id[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.850 323.915 49.130 327.915 ;
    END
  END arbitration_id[16]
  PIN arbitration_id[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 51.150 323.915 51.430 327.915 ;
    END
  END arbitration_id[17]
  PIN arbitration_id[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 53.450 323.915 53.730 327.915 ;
    END
  END arbitration_id[18]
  PIN arbitration_id[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 55.750 323.915 56.030 327.915 ;
    END
  END arbitration_id[19]
  PIN arbitration_id[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 14.350 323.915 14.630 327.915 ;
    END
  END arbitration_id[1]
  PIN arbitration_id[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 323.915 58.330 327.915 ;
    END
  END arbitration_id[20]
  PIN arbitration_id[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 60.350 323.915 60.630 327.915 ;
    END
  END arbitration_id[21]
  PIN arbitration_id[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 62.650 323.915 62.930 327.915 ;
    END
  END arbitration_id[22]
  PIN arbitration_id[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.950 323.915 65.230 327.915 ;
    END
  END arbitration_id[23]
  PIN arbitration_id[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.250 323.915 67.530 327.915 ;
    END
  END arbitration_id[24]
  PIN arbitration_id[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 69.550 323.915 69.830 327.915 ;
    END
  END arbitration_id[25]
  PIN arbitration_id[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 71.850 323.915 72.130 327.915 ;
    END
  END arbitration_id[26]
  PIN arbitration_id[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 74.150 323.915 74.430 327.915 ;
    END
  END arbitration_id[27]
  PIN arbitration_id[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 76.450 323.915 76.730 327.915 ;
    END
  END arbitration_id[28]
  PIN arbitration_id[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 78.750 323.915 79.030 327.915 ;
    END
  END arbitration_id[29]
  PIN arbitration_id[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.650 323.915 16.930 327.915 ;
    END
  END arbitration_id[2]
  PIN arbitration_id[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 81.050 323.915 81.330 327.915 ;
    END
  END arbitration_id[30]
  PIN arbitration_id[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.350 323.915 83.630 327.915 ;
    END
  END arbitration_id[31]
  PIN arbitration_id[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 85.650 323.915 85.930 327.915 ;
    END
  END arbitration_id[32]
  PIN arbitration_id[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.950 323.915 88.230 327.915 ;
    END
  END arbitration_id[33]
  PIN arbitration_id[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 323.915 90.530 327.915 ;
    END
  END arbitration_id[34]
  PIN arbitration_id[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 92.550 323.915 92.830 327.915 ;
    END
  END arbitration_id[35]
  PIN arbitration_id[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 94.850 323.915 95.130 327.915 ;
    END
  END arbitration_id[36]
  PIN arbitration_id[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 97.150 323.915 97.430 327.915 ;
    END
  END arbitration_id[37]
  PIN arbitration_id[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.450 323.915 99.730 327.915 ;
    END
  END arbitration_id[38]
  PIN arbitration_id[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 101.750 323.915 102.030 327.915 ;
    END
  END arbitration_id[39]
  PIN arbitration_id[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 18.950 323.915 19.230 327.915 ;
    END
  END arbitration_id[3]
  PIN arbitration_id[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 104.050 323.915 104.330 327.915 ;
    END
  END arbitration_id[40]
  PIN arbitration_id[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 323.915 106.630 327.915 ;
    END
  END arbitration_id[41]
  PIN arbitration_id[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 108.650 323.915 108.930 327.915 ;
    END
  END arbitration_id[42]
  PIN arbitration_id[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 110.950 323.915 111.230 327.915 ;
    END
  END arbitration_id[43]
  PIN arbitration_id[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 113.250 323.915 113.530 327.915 ;
    END
  END arbitration_id[44]
  PIN arbitration_id[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 115.550 323.915 115.830 327.915 ;
    END
  END arbitration_id[45]
  PIN arbitration_id[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 117.850 323.915 118.130 327.915 ;
    END
  END arbitration_id[46]
  PIN arbitration_id[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 120.150 323.915 120.430 327.915 ;
    END
  END arbitration_id[47]
  PIN arbitration_id[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 323.915 122.730 327.915 ;
    END
  END arbitration_id[48]
  PIN arbitration_id[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 124.750 323.915 125.030 327.915 ;
    END
  END arbitration_id[49]
  PIN arbitration_id[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 21.250 323.915 21.530 327.915 ;
    END
  END arbitration_id[4]
  PIN arbitration_id[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 127.050 323.915 127.330 327.915 ;
    END
  END arbitration_id[50]
  PIN arbitration_id[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 129.350 323.915 129.630 327.915 ;
    END
  END arbitration_id[51]
  PIN arbitration_id[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 131.650 323.915 131.930 327.915 ;
    END
  END arbitration_id[52]
  PIN arbitration_id[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 133.950 323.915 134.230 327.915 ;
    END
  END arbitration_id[53]
  PIN arbitration_id[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 136.250 323.915 136.530 327.915 ;
    END
  END arbitration_id[54]
  PIN arbitration_id[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 323.915 138.830 327.915 ;
    END
  END arbitration_id[55]
  PIN arbitration_id[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 140.850 323.915 141.130 327.915 ;
    END
  END arbitration_id[56]
  PIN arbitration_id[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 143.150 323.915 143.430 327.915 ;
    END
  END arbitration_id[57]
  PIN arbitration_id[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 145.450 323.915 145.730 327.915 ;
    END
  END arbitration_id[58]
  PIN arbitration_id[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 147.750 323.915 148.030 327.915 ;
    END
  END arbitration_id[59]
  PIN arbitration_id[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 23.550 323.915 23.830 327.915 ;
    END
  END arbitration_id[5]
  PIN arbitration_id[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 150.050 323.915 150.330 327.915 ;
    END
  END arbitration_id[60]
  PIN arbitration_id[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 152.350 323.915 152.630 327.915 ;
    END
  END arbitration_id[61]
  PIN arbitration_id[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 323.915 154.930 327.915 ;
    END
  END arbitration_id[62]
  PIN arbitration_id[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 156.950 323.915 157.230 327.915 ;
    END
  END arbitration_id[63]
  PIN arbitration_id[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 323.915 26.130 327.915 ;
    END
  END arbitration_id[6]
  PIN arbitration_id[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 28.150 323.915 28.430 327.915 ;
    END
  END arbitration_id[7]
  PIN arbitration_id[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 30.450 323.915 30.730 327.915 ;
    END
  END arbitration_id[8]
  PIN arbitration_id[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.750 323.915 33.030 327.915 ;
    END
  END arbitration_id[9]
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 79.210 0.000 79.490 4.000 ;
    END
  END clk
  PIN data_field[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 29.960 317.195 30.560 ;
    END
  END data_field[0]
  PIN data_field[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 70.760 317.195 71.360 ;
    END
  END data_field[10]
  PIN data_field[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 74.840 317.195 75.440 ;
    END
  END data_field[11]
  PIN data_field[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 78.920 317.195 79.520 ;
    END
  END data_field[12]
  PIN data_field[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 83.000 317.195 83.600 ;
    END
  END data_field[13]
  PIN data_field[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 87.080 317.195 87.680 ;
    END
  END data_field[14]
  PIN data_field[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 91.160 317.195 91.760 ;
    END
  END data_field[15]
  PIN data_field[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 95.240 317.195 95.840 ;
    END
  END data_field[16]
  PIN data_field[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 99.320 317.195 99.920 ;
    END
  END data_field[17]
  PIN data_field[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 103.400 317.195 104.000 ;
    END
  END data_field[18]
  PIN data_field[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 107.480 317.195 108.080 ;
    END
  END data_field[19]
  PIN data_field[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 34.040 317.195 34.640 ;
    END
  END data_field[1]
  PIN data_field[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 111.560 317.195 112.160 ;
    END
  END data_field[20]
  PIN data_field[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 115.640 317.195 116.240 ;
    END
  END data_field[21]
  PIN data_field[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 119.720 317.195 120.320 ;
    END
  END data_field[22]
  PIN data_field[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 123.800 317.195 124.400 ;
    END
  END data_field[23]
  PIN data_field[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 127.880 317.195 128.480 ;
    END
  END data_field[24]
  PIN data_field[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 131.960 317.195 132.560 ;
    END
  END data_field[25]
  PIN data_field[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 136.040 317.195 136.640 ;
    END
  END data_field[26]
  PIN data_field[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 140.120 317.195 140.720 ;
    END
  END data_field[27]
  PIN data_field[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 144.200 317.195 144.800 ;
    END
  END data_field[28]
  PIN data_field[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 148.280 317.195 148.880 ;
    END
  END data_field[29]
  PIN data_field[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 38.120 317.195 38.720 ;
    END
  END data_field[2]
  PIN data_field[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 152.360 317.195 152.960 ;
    END
  END data_field[30]
  PIN data_field[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 156.440 317.195 157.040 ;
    END
  END data_field[31]
  PIN data_field[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 160.520 317.195 161.120 ;
    END
  END data_field[32]
  PIN data_field[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 164.600 317.195 165.200 ;
    END
  END data_field[33]
  PIN data_field[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 168.680 317.195 169.280 ;
    END
  END data_field[34]
  PIN data_field[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 172.760 317.195 173.360 ;
    END
  END data_field[35]
  PIN data_field[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 176.840 317.195 177.440 ;
    END
  END data_field[36]
  PIN data_field[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 180.920 317.195 181.520 ;
    END
  END data_field[37]
  PIN data_field[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 185.000 317.195 185.600 ;
    END
  END data_field[38]
  PIN data_field[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 189.080 317.195 189.680 ;
    END
  END data_field[39]
  PIN data_field[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 42.200 317.195 42.800 ;
    END
  END data_field[3]
  PIN data_field[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 193.160 317.195 193.760 ;
    END
  END data_field[40]
  PIN data_field[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 197.240 317.195 197.840 ;
    END
  END data_field[41]
  PIN data_field[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 201.320 317.195 201.920 ;
    END
  END data_field[42]
  PIN data_field[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 205.400 317.195 206.000 ;
    END
  END data_field[43]
  PIN data_field[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 209.480 317.195 210.080 ;
    END
  END data_field[44]
  PIN data_field[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 213.560 317.195 214.160 ;
    END
  END data_field[45]
  PIN data_field[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 217.640 317.195 218.240 ;
    END
  END data_field[46]
  PIN data_field[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 221.720 317.195 222.320 ;
    END
  END data_field[47]
  PIN data_field[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 225.800 317.195 226.400 ;
    END
  END data_field[48]
  PIN data_field[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 229.880 317.195 230.480 ;
    END
  END data_field[49]
  PIN data_field[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 46.280 317.195 46.880 ;
    END
  END data_field[4]
  PIN data_field[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 233.960 317.195 234.560 ;
    END
  END data_field[50]
  PIN data_field[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 238.040 317.195 238.640 ;
    END
  END data_field[51]
  PIN data_field[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 242.120 317.195 242.720 ;
    END
  END data_field[52]
  PIN data_field[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 246.200 317.195 246.800 ;
    END
  END data_field[53]
  PIN data_field[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 250.280 317.195 250.880 ;
    END
  END data_field[54]
  PIN data_field[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 254.360 317.195 254.960 ;
    END
  END data_field[55]
  PIN data_field[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 258.440 317.195 259.040 ;
    END
  END data_field[56]
  PIN data_field[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 262.520 317.195 263.120 ;
    END
  END data_field[57]
  PIN data_field[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 266.600 317.195 267.200 ;
    END
  END data_field[58]
  PIN data_field[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 270.680 317.195 271.280 ;
    END
  END data_field[59]
  PIN data_field[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 50.360 317.195 50.960 ;
    END
  END data_field[5]
  PIN data_field[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 274.760 317.195 275.360 ;
    END
  END data_field[60]
  PIN data_field[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 278.840 317.195 279.440 ;
    END
  END data_field[61]
  PIN data_field[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 282.920 317.195 283.520 ;
    END
  END data_field[62]
  PIN data_field[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 287.000 317.195 287.600 ;
    END
  END data_field[63]
  PIN data_field[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 54.440 317.195 55.040 ;
    END
  END data_field[6]
  PIN data_field[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 58.520 317.195 59.120 ;
    END
  END data_field[7]
  PIN data_field[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 62.600 317.195 63.200 ;
    END
  END data_field[8]
  PIN data_field[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 313.195 66.680 317.195 67.280 ;
    END
  END data_field[9]
  PIN feature_valid
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met3 ;
        RECT 313.195 291.080 317.195 291.680 ;
    END
  END feature_valid
  PIN frame_id_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.000 4.000 117.600 ;
    END
  END frame_id_out[0]
  PIN frame_id_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 163.240 4.000 163.840 ;
    END
  END frame_id_out[1]
  PIN frame_id_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 209.480 4.000 210.080 ;
    END
  END frame_id_out[2]
  PIN frame_id_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END frame_id_out[3]
  PIN frame_id_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END frame_id_out[4]
  PIN prediction_out
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.760 4.000 71.360 ;
    END
  END prediction_out
  PIN prediction_valid
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END prediction_valid
  PIN ready_for_next
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.782000 ;
    PORT
      LAYER met3 ;
        RECT 313.195 295.160 317.195 295.760 ;
    END
  END ready_for_next
  PIN rst_n
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.990000 ;
    ANTENNADIFFAREA 0.434700 ;
    PORT
      LAYER met2 ;
        RECT 237.450 0.000 237.730 4.000 ;
    END
  END rst_n
  PIN timestamp[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 159.250 323.915 159.530 327.915 ;
    END
  END timestamp[0]
  PIN timestamp[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 182.250 323.915 182.530 327.915 ;
    END
  END timestamp[10]
  PIN timestamp[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 184.550 323.915 184.830 327.915 ;
    END
  END timestamp[11]
  PIN timestamp[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 186.850 323.915 187.130 327.915 ;
    END
  END timestamp[12]
  PIN timestamp[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 189.150 323.915 189.430 327.915 ;
    END
  END timestamp[13]
  PIN timestamp[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 191.450 323.915 191.730 327.915 ;
    END
  END timestamp[14]
  PIN timestamp[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.750 323.915 194.030 327.915 ;
    END
  END timestamp[15]
  PIN timestamp[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.050 323.915 196.330 327.915 ;
    END
  END timestamp[16]
  PIN timestamp[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 198.350 323.915 198.630 327.915 ;
    END
  END timestamp[17]
  PIN timestamp[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 200.650 323.915 200.930 327.915 ;
    END
  END timestamp[18]
  PIN timestamp[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 323.915 203.230 327.915 ;
    END
  END timestamp[19]
  PIN timestamp[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.550 323.915 161.830 327.915 ;
    END
  END timestamp[1]
  PIN timestamp[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 205.250 323.915 205.530 327.915 ;
    END
  END timestamp[20]
  PIN timestamp[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 207.550 323.915 207.830 327.915 ;
    END
  END timestamp[21]
  PIN timestamp[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 209.850 323.915 210.130 327.915 ;
    END
  END timestamp[22]
  PIN timestamp[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.150 323.915 212.430 327.915 ;
    END
  END timestamp[23]
  PIN timestamp[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 214.450 323.915 214.730 327.915 ;
    END
  END timestamp[24]
  PIN timestamp[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 216.750 323.915 217.030 327.915 ;
    END
  END timestamp[25]
  PIN timestamp[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 323.915 219.330 327.915 ;
    END
  END timestamp[26]
  PIN timestamp[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 221.350 323.915 221.630 327.915 ;
    END
  END timestamp[27]
  PIN timestamp[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 223.650 323.915 223.930 327.915 ;
    END
  END timestamp[28]
  PIN timestamp[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.950 323.915 226.230 327.915 ;
    END
  END timestamp[29]
  PIN timestamp[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 163.850 323.915 164.130 327.915 ;
    END
  END timestamp[2]
  PIN timestamp[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.250 323.915 228.530 327.915 ;
    END
  END timestamp[30]
  PIN timestamp[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 230.550 323.915 230.830 327.915 ;
    END
  END timestamp[31]
  PIN timestamp[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 232.850 323.915 233.130 327.915 ;
    END
  END timestamp[32]
  PIN timestamp[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 323.915 235.430 327.915 ;
    END
  END timestamp[33]
  PIN timestamp[34]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 237.450 323.915 237.730 327.915 ;
    END
  END timestamp[34]
  PIN timestamp[35]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 239.750 323.915 240.030 327.915 ;
    END
  END timestamp[35]
  PIN timestamp[36]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 242.050 323.915 242.330 327.915 ;
    END
  END timestamp[36]
  PIN timestamp[37]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.350 323.915 244.630 327.915 ;
    END
  END timestamp[37]
  PIN timestamp[38]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 246.650 323.915 246.930 327.915 ;
    END
  END timestamp[38]
  PIN timestamp[39]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.950 323.915 249.230 327.915 ;
    END
  END timestamp[39]
  PIN timestamp[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 166.150 323.915 166.430 327.915 ;
    END
  END timestamp[3]
  PIN timestamp[40]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 323.915 251.530 327.915 ;
    END
  END timestamp[40]
  PIN timestamp[41]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 253.550 323.915 253.830 327.915 ;
    END
  END timestamp[41]
  PIN timestamp[42]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 255.850 323.915 256.130 327.915 ;
    END
  END timestamp[42]
  PIN timestamp[43]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 258.150 323.915 258.430 327.915 ;
    END
  END timestamp[43]
  PIN timestamp[44]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.450 323.915 260.730 327.915 ;
    END
  END timestamp[44]
  PIN timestamp[45]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 262.750 323.915 263.030 327.915 ;
    END
  END timestamp[45]
  PIN timestamp[46]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 265.050 323.915 265.330 327.915 ;
    END
  END timestamp[46]
  PIN timestamp[47]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 323.915 267.630 327.915 ;
    END
  END timestamp[47]
  PIN timestamp[48]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 269.650 323.915 269.930 327.915 ;
    END
  END timestamp[48]
  PIN timestamp[49]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 271.950 323.915 272.230 327.915 ;
    END
  END timestamp[49]
  PIN timestamp[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 168.450 323.915 168.730 327.915 ;
    END
  END timestamp[4]
  PIN timestamp[50]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 274.250 323.915 274.530 327.915 ;
    END
  END timestamp[50]
  PIN timestamp[51]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 276.550 323.915 276.830 327.915 ;
    END
  END timestamp[51]
  PIN timestamp[52]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 278.850 323.915 279.130 327.915 ;
    END
  END timestamp[52]
  PIN timestamp[53]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 281.150 323.915 281.430 327.915 ;
    END
  END timestamp[53]
  PIN timestamp[54]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 323.915 283.730 327.915 ;
    END
  END timestamp[54]
  PIN timestamp[55]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 285.750 323.915 286.030 327.915 ;
    END
  END timestamp[55]
  PIN timestamp[56]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 288.050 323.915 288.330 327.915 ;
    END
  END timestamp[56]
  PIN timestamp[57]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 290.350 323.915 290.630 327.915 ;
    END
  END timestamp[57]
  PIN timestamp[58]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 292.650 323.915 292.930 327.915 ;
    END
  END timestamp[58]
  PIN timestamp[59]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 294.950 323.915 295.230 327.915 ;
    END
  END timestamp[59]
  PIN timestamp[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 323.915 171.030 327.915 ;
    END
  END timestamp[5]
  PIN timestamp[60]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 297.250 323.915 297.530 327.915 ;
    END
  END timestamp[60]
  PIN timestamp[61]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 323.915 299.830 327.915 ;
    END
  END timestamp[61]
  PIN timestamp[62]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 301.850 323.915 302.130 327.915 ;
    END
  END timestamp[62]
  PIN timestamp[63]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 304.150 323.915 304.430 327.915 ;
    END
  END timestamp[63]
  PIN timestamp[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.050 323.915 173.330 327.915 ;
    END
  END timestamp[6]
  PIN timestamp[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 175.350 323.915 175.630 327.915 ;
    END
  END timestamp[7]
  PIN timestamp[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.650 323.915 177.930 327.915 ;
    END
  END timestamp[8]
  PIN timestamp[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 179.950 323.915 180.230 327.915 ;
    END
  END timestamp[9]
  OBS
      LAYER nwell ;
        RECT 5.330 10.795 311.610 315.605 ;
      LAYER li1 ;
        RECT 5.520 10.795 311.420 315.605 ;
      LAYER met1 ;
        RECT 4.210 10.640 312.730 315.760 ;
      LAYER met2 ;
        RECT 4.230 4.280 312.710 315.705 ;
        RECT 4.230 4.000 78.930 4.280 ;
        RECT 79.770 4.000 237.170 4.280 ;
        RECT 238.010 4.000 312.710 4.280 ;
      LAYER met3 ;
        RECT 3.990 302.960 313.195 315.685 ;
        RECT 4.400 301.560 313.195 302.960 ;
        RECT 3.990 296.160 313.195 301.560 ;
        RECT 3.990 294.760 312.795 296.160 ;
        RECT 3.990 292.080 313.195 294.760 ;
        RECT 3.990 290.680 312.795 292.080 ;
        RECT 3.990 288.000 313.195 290.680 ;
        RECT 3.990 286.600 312.795 288.000 ;
        RECT 3.990 283.920 313.195 286.600 ;
        RECT 3.990 282.520 312.795 283.920 ;
        RECT 3.990 279.840 313.195 282.520 ;
        RECT 3.990 278.440 312.795 279.840 ;
        RECT 3.990 275.760 313.195 278.440 ;
        RECT 3.990 274.360 312.795 275.760 ;
        RECT 3.990 271.680 313.195 274.360 ;
        RECT 3.990 270.280 312.795 271.680 ;
        RECT 3.990 267.600 313.195 270.280 ;
        RECT 3.990 266.200 312.795 267.600 ;
        RECT 3.990 263.520 313.195 266.200 ;
        RECT 3.990 262.120 312.795 263.520 ;
        RECT 3.990 259.440 313.195 262.120 ;
        RECT 3.990 258.040 312.795 259.440 ;
        RECT 3.990 256.720 313.195 258.040 ;
        RECT 4.400 255.360 313.195 256.720 ;
        RECT 4.400 255.320 312.795 255.360 ;
        RECT 3.990 253.960 312.795 255.320 ;
        RECT 3.990 251.280 313.195 253.960 ;
        RECT 3.990 249.880 312.795 251.280 ;
        RECT 3.990 247.200 313.195 249.880 ;
        RECT 3.990 245.800 312.795 247.200 ;
        RECT 3.990 243.120 313.195 245.800 ;
        RECT 3.990 241.720 312.795 243.120 ;
        RECT 3.990 239.040 313.195 241.720 ;
        RECT 3.990 237.640 312.795 239.040 ;
        RECT 3.990 234.960 313.195 237.640 ;
        RECT 3.990 233.560 312.795 234.960 ;
        RECT 3.990 230.880 313.195 233.560 ;
        RECT 3.990 229.480 312.795 230.880 ;
        RECT 3.990 226.800 313.195 229.480 ;
        RECT 3.990 225.400 312.795 226.800 ;
        RECT 3.990 222.720 313.195 225.400 ;
        RECT 3.990 221.320 312.795 222.720 ;
        RECT 3.990 218.640 313.195 221.320 ;
        RECT 3.990 217.240 312.795 218.640 ;
        RECT 3.990 214.560 313.195 217.240 ;
        RECT 3.990 213.160 312.795 214.560 ;
        RECT 3.990 210.480 313.195 213.160 ;
        RECT 4.400 209.080 312.795 210.480 ;
        RECT 3.990 206.400 313.195 209.080 ;
        RECT 3.990 205.000 312.795 206.400 ;
        RECT 3.990 202.320 313.195 205.000 ;
        RECT 3.990 200.920 312.795 202.320 ;
        RECT 3.990 198.240 313.195 200.920 ;
        RECT 3.990 196.840 312.795 198.240 ;
        RECT 3.990 194.160 313.195 196.840 ;
        RECT 3.990 192.760 312.795 194.160 ;
        RECT 3.990 190.080 313.195 192.760 ;
        RECT 3.990 188.680 312.795 190.080 ;
        RECT 3.990 186.000 313.195 188.680 ;
        RECT 3.990 184.600 312.795 186.000 ;
        RECT 3.990 181.920 313.195 184.600 ;
        RECT 3.990 180.520 312.795 181.920 ;
        RECT 3.990 177.840 313.195 180.520 ;
        RECT 3.990 176.440 312.795 177.840 ;
        RECT 3.990 173.760 313.195 176.440 ;
        RECT 3.990 172.360 312.795 173.760 ;
        RECT 3.990 169.680 313.195 172.360 ;
        RECT 3.990 168.280 312.795 169.680 ;
        RECT 3.990 165.600 313.195 168.280 ;
        RECT 3.990 164.240 312.795 165.600 ;
        RECT 4.400 164.200 312.795 164.240 ;
        RECT 4.400 162.840 313.195 164.200 ;
        RECT 3.990 161.520 313.195 162.840 ;
        RECT 3.990 160.120 312.795 161.520 ;
        RECT 3.990 157.440 313.195 160.120 ;
        RECT 3.990 156.040 312.795 157.440 ;
        RECT 3.990 153.360 313.195 156.040 ;
        RECT 3.990 151.960 312.795 153.360 ;
        RECT 3.990 149.280 313.195 151.960 ;
        RECT 3.990 147.880 312.795 149.280 ;
        RECT 3.990 145.200 313.195 147.880 ;
        RECT 3.990 143.800 312.795 145.200 ;
        RECT 3.990 141.120 313.195 143.800 ;
        RECT 3.990 139.720 312.795 141.120 ;
        RECT 3.990 137.040 313.195 139.720 ;
        RECT 3.990 135.640 312.795 137.040 ;
        RECT 3.990 132.960 313.195 135.640 ;
        RECT 3.990 131.560 312.795 132.960 ;
        RECT 3.990 128.880 313.195 131.560 ;
        RECT 3.990 127.480 312.795 128.880 ;
        RECT 3.990 124.800 313.195 127.480 ;
        RECT 3.990 123.400 312.795 124.800 ;
        RECT 3.990 120.720 313.195 123.400 ;
        RECT 3.990 119.320 312.795 120.720 ;
        RECT 3.990 118.000 313.195 119.320 ;
        RECT 4.400 116.640 313.195 118.000 ;
        RECT 4.400 116.600 312.795 116.640 ;
        RECT 3.990 115.240 312.795 116.600 ;
        RECT 3.990 112.560 313.195 115.240 ;
        RECT 3.990 111.160 312.795 112.560 ;
        RECT 3.990 108.480 313.195 111.160 ;
        RECT 3.990 107.080 312.795 108.480 ;
        RECT 3.990 104.400 313.195 107.080 ;
        RECT 3.990 103.000 312.795 104.400 ;
        RECT 3.990 100.320 313.195 103.000 ;
        RECT 3.990 98.920 312.795 100.320 ;
        RECT 3.990 96.240 313.195 98.920 ;
        RECT 3.990 94.840 312.795 96.240 ;
        RECT 3.990 92.160 313.195 94.840 ;
        RECT 3.990 90.760 312.795 92.160 ;
        RECT 3.990 88.080 313.195 90.760 ;
        RECT 3.990 86.680 312.795 88.080 ;
        RECT 3.990 84.000 313.195 86.680 ;
        RECT 3.990 82.600 312.795 84.000 ;
        RECT 3.990 79.920 313.195 82.600 ;
        RECT 3.990 78.520 312.795 79.920 ;
        RECT 3.990 75.840 313.195 78.520 ;
        RECT 3.990 74.440 312.795 75.840 ;
        RECT 3.990 71.760 313.195 74.440 ;
        RECT 4.400 70.360 312.795 71.760 ;
        RECT 3.990 67.680 313.195 70.360 ;
        RECT 3.990 66.280 312.795 67.680 ;
        RECT 3.990 63.600 313.195 66.280 ;
        RECT 3.990 62.200 312.795 63.600 ;
        RECT 3.990 59.520 313.195 62.200 ;
        RECT 3.990 58.120 312.795 59.520 ;
        RECT 3.990 55.440 313.195 58.120 ;
        RECT 3.990 54.040 312.795 55.440 ;
        RECT 3.990 51.360 313.195 54.040 ;
        RECT 3.990 49.960 312.795 51.360 ;
        RECT 3.990 47.280 313.195 49.960 ;
        RECT 3.990 45.880 312.795 47.280 ;
        RECT 3.990 43.200 313.195 45.880 ;
        RECT 3.990 41.800 312.795 43.200 ;
        RECT 3.990 39.120 313.195 41.800 ;
        RECT 3.990 37.720 312.795 39.120 ;
        RECT 3.990 35.040 313.195 37.720 ;
        RECT 3.990 33.640 312.795 35.040 ;
        RECT 3.990 30.960 313.195 33.640 ;
        RECT 3.990 29.560 312.795 30.960 ;
        RECT 3.990 25.520 313.195 29.560 ;
        RECT 4.400 24.120 313.195 25.520 ;
        RECT 3.990 10.715 313.195 24.120 ;
      LAYER met4 ;
        RECT 17.775 17.175 38.620 303.785 ;
        RECT 42.420 17.175 43.320 303.785 ;
        RECT 47.120 17.175 68.620 303.785 ;
        RECT 72.420 17.175 73.320 303.785 ;
        RECT 77.120 17.175 98.620 303.785 ;
        RECT 102.420 17.175 103.320 303.785 ;
        RECT 107.120 17.175 128.620 303.785 ;
        RECT 132.420 17.175 133.320 303.785 ;
        RECT 137.120 17.175 158.620 303.785 ;
        RECT 162.420 17.175 163.320 303.785 ;
        RECT 167.120 17.175 188.620 303.785 ;
        RECT 192.420 17.175 193.320 303.785 ;
        RECT 197.120 17.175 218.620 303.785 ;
        RECT 222.420 17.175 223.320 303.785 ;
        RECT 227.120 17.175 248.620 303.785 ;
        RECT 252.420 17.175 253.320 303.785 ;
        RECT 257.120 17.175 278.620 303.785 ;
        RECT 282.420 17.175 283.320 303.785 ;
        RECT 287.120 17.175 289.505 303.785 ;
  END
END Random_forest_top_ver2
END LIBRARY

