module tree_rom_9 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000041D8EC33900000000010CC3;
    rom[1] = 120'h001140681000000000000020033;
    rom[2] = 120'h002300000000000000000000001;
    rom[3] = 120'h003041D8EC335000000000405B3;
    rom[4] = 120'h004A43D46E4A6000000000503C3;
    rom[5] = 120'h005A4170180BC000000000601D3;
    rom[6] = 120'h006A41385AA8800000000070143;
    rom[7] = 120'h007A40EFFD400000000000800F3;
    rom[8] = 120'h008A400400000000000000900C3;
    rom[9] = 120'h009A3FF800000000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000000;
    rom[12] = 120'h00C1407348000000000000D00E3;
    rom[13] = 120'h00D300000000000000000000001;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00F1407F8800000000000100133;
    rom[16] = 120'h010A4134EA94800000000110123;
    rom[17] = 120'h011300000000000000000000000;
    rom[18] = 120'h012300000000000000000000000;
    rom[19] = 120'h013300000000000000000000001;
    rom[20] = 120'h0141408A58000000000001501C3;
    rom[21] = 120'h0151408A3C00000000000160193;
    rom[22] = 120'h01614079E000000000000170183;
    rom[23] = 120'h017300000000000000000000001;
    rom[24] = 120'h018300000000000000000000001;
    rom[25] = 120'h019A415794C6E000000001A01B3;
    rom[26] = 120'h01A300000000000000000000001;
    rom[27] = 120'h01B300000000000000000000000;
    rom[28] = 120'h01C300000000000000000000001;
    rom[29] = 120'h01DA435FFC444000000001E02D3;
    rom[30] = 120'h01E1407E18000000000001F0263;
    rom[31] = 120'h01FA41EF934BC00000000200233;
    rom[32] = 120'h0201406E1000000000000210223;
    rom[33] = 120'h021300000000000000000000001;
    rom[34] = 120'h022300000000000000000000000;
    rom[35] = 120'h023140783800000000000240253;
    rom[36] = 120'h024300000000000000000000000;
    rom[37] = 120'h025300000000000000000000000;
    rom[38] = 120'h0261408A54000000000002702A3;
    rom[39] = 120'h027140861400000000000280293;
    rom[40] = 120'h028300000000000000000000001;
    rom[41] = 120'h029300000000000000000000000;
    rom[42] = 120'h02AA426C1C6AE000000002B02C3;
    rom[43] = 120'h02B300000000000000000000001;
    rom[44] = 120'h02C300000000000000000000001;
    rom[45] = 120'h02D1407F58000000000002E0353;
    rom[46] = 120'h02E1406930000000000002F0323;
    rom[47] = 120'h02FA43CA7D45B00000000300313;
    rom[48] = 120'h030300000000000000000000000;
    rom[49] = 120'h031300000000000000000000001;
    rom[50] = 120'h032140790800000000000330343;
    rom[51] = 120'h033300000000000000000000001;
    rom[52] = 120'h034300000000000000000000000;
    rom[53] = 120'h035A43A007F9500000000360393;
    rom[54] = 120'h0361408F8C00000000000370383;
    rom[55] = 120'h037300000000000000000000000;
    rom[56] = 120'h038300000000000000000000001;
    rom[57] = 120'h03914094AA000000000003A03B3;
    rom[58] = 120'h03A300000000000000000000001;
    rom[59] = 120'h03B300000000000000000000001;
    rom[60] = 120'h03C1407F18000000000003D0523;
    rom[61] = 120'h03DA43DEDB482000000003E0453;
    rom[62] = 120'h03EA43D5BB4E3000000003F0403;
    rom[63] = 120'h03F300000000000000000000001;
    rom[64] = 120'h040A43D5C16F300000000410423;
    rom[65] = 120'h041300000000000000000000000;
    rom[66] = 120'h042A43D5FF24400000000430443;
    rom[67] = 120'h043300000000000000000000001;
    rom[68] = 120'h044300000000000000000000001;
    rom[69] = 120'h045A43EA38339000000004604D3;
    rom[70] = 120'h0461407980000000000004704A3;
    rom[71] = 120'h0471406F3000000000000480493;
    rom[72] = 120'h048300000000000000000000000;
    rom[73] = 120'h049300000000000000000000001;
    rom[74] = 120'h04A14079D8000000000004B04C3;
    rom[75] = 120'h04B300000000000000000000000;
    rom[76] = 120'h04C300000000000000000000001;
    rom[77] = 120'h04D1407988000000000004E04F3;
    rom[78] = 120'h04E300000000000000000000001;
    rom[79] = 120'h04FA43EAF9AD900000000500513;
    rom[80] = 120'h050300000000000000000000001;
    rom[81] = 120'h051300000000000000000000001;
    rom[82] = 120'h0521408F6C000000000005305A3;
    rom[83] = 120'h0531408F6400000000000540553;
    rom[84] = 120'h054300000000000000000000001;
    rom[85] = 120'h055A43DF0C73100000000560573;
    rom[86] = 120'h056300000000000000000000001;
    rom[87] = 120'h057A43E316E8A00000000580593;
    rom[88] = 120'h058300000000000000000000000;
    rom[89] = 120'h059300000000000000000000001;
    rom[90] = 120'h05A300000000000000000000001;
    rom[91] = 120'h05B1407E58000000000005C0953;
    rom[92] = 120'h05CA40EFE0F00000000005D07A3;
    rom[93] = 120'h05D1407338000000000005E06B3;
    rom[94] = 120'h05E041D8EC337000000005F0663;
    rom[95] = 120'h05F14068B000000000000600633;
    rom[96] = 120'h060140689000000000000610623;
    rom[97] = 120'h061300000000000000000000000;
    rom[98] = 120'h062300000000000000000000000;
    rom[99] = 120'h063A40CED280000000000640653;
    rom[100] = 120'h064300000000000000000000001;
    rom[101] = 120'h065300000000000000000000000;
    rom[102] = 120'h0661406DF000000000000670683;
    rom[103] = 120'h067300000000000000000000001;
    rom[104] = 120'h068A405040000000000006906A3;
    rom[105] = 120'h069300000000000000000000000;
    rom[106] = 120'h06A300000000000000000000001;
    rom[107] = 120'h06B14077E8000000000006C0733;
    rom[108] = 120'h06CA40A6B6000000000006D0703;
    rom[109] = 120'h06D1407388000000000006E06F3;
    rom[110] = 120'h06E300000000000000000000000;
    rom[111] = 120'h06F300000000000000000000001;
    rom[112] = 120'h070140736800000000000710723;
    rom[113] = 120'h071300000000000000000000000;
    rom[114] = 120'h072300000000000000000000001;
    rom[115] = 120'h073041D8EC33700000000740773;
    rom[116] = 120'h074A404FC000000000000750763;
    rom[117] = 120'h075300000000000000000000000;
    rom[118] = 120'h076300000000000000000000001;
    rom[119] = 120'h0771407CE000000000000780793;
    rom[120] = 120'h078300000000000000000000000;
    rom[121] = 120'h079300000000000000000000001;
    rom[122] = 120'h07A041D8EC337000000007B0883;
    rom[123] = 120'h07BA43D3FFF05000000007C0833;
    rom[124] = 120'h07C14077C8000000000007D0803;
    rom[125] = 120'h07D1406F30000000000007E07F3;
    rom[126] = 120'h07E300000000000000000000000;
    rom[127] = 120'h07F300000000000000000000001;
    rom[128] = 120'h0801407E0800000000000810823;
    rom[129] = 120'h081300000000000000000000000;
    rom[130] = 120'h082300000000000000000000000;
    rom[131] = 120'h083140798800000000000840853;
    rom[132] = 120'h084300000000000000000000001;
    rom[133] = 120'h085A43DFFABFC00000000860873;
    rom[134] = 120'h086300000000000000000000001;
    rom[135] = 120'h087300000000000000000000000;
    rom[136] = 120'h088A43E20BB1000000000890903;
    rom[137] = 120'h089A436080074000000008A08D3;
    rom[138] = 120'h08A1407838000000000008B08C3;
    rom[139] = 120'h08B300000000000000000000000;
    rom[140] = 120'h08C300000000000000000000000;
    rom[141] = 120'h08DA43C21300C000000008E08F3;
    rom[142] = 120'h08E300000000000000000000000;
    rom[143] = 120'h08F300000000000000000000000;
    rom[144] = 120'h090140798000000000000910923;
    rom[145] = 120'h091300000000000000000000001;
    rom[146] = 120'h092A43EA163C600000000930943;
    rom[147] = 120'h093300000000000000000000000;
    rom[148] = 120'h094300000000000000000000001;
    rom[149] = 120'h0951408E8C00000000000960AD3;
    rom[150] = 120'h096A3FE000000000000009709E3;
    rom[151] = 120'h097041D8EC337000000009809D3;
    rom[152] = 120'h09814088D4000000000009909C3;
    rom[153] = 120'h0991408104000000000009A09B3;
    rom[154] = 120'h09A300000000000000000000000;
    rom[155] = 120'h09B300000000000000000000001;
    rom[156] = 120'h09C300000000000000000000000;
    rom[157] = 120'h09D300000000000000000000000;
    rom[158] = 120'h09E041D8EC337000000009F0A63;
    rom[159] = 120'h09F1408E0400000000000A00A33;
    rom[160] = 120'h0A01408A5400000000000A10A23;
    rom[161] = 120'h0A1300000000000000000000001;
    rom[162] = 120'h0A2300000000000000000000001;
    rom[163] = 120'h0A3A4374B000000000000A40A53;
    rom[164] = 120'h0A4300000000000000000000001;
    rom[165] = 120'h0A5300000000000000000000000;
    rom[166] = 120'h0A6A42A27543C00000000A70AA3;
    rom[167] = 120'h0A7A416BF44EF00000000A80A93;
    rom[168] = 120'h0A8300000000000000000000001;
    rom[169] = 120'h0A9300000000000000000000000;
    rom[170] = 120'h0AAA43AE3600300000000AB0AC3;
    rom[171] = 120'h0AB300000000000000000000001;
    rom[172] = 120'h0AC300000000000000000000000;
    rom[173] = 120'h0AD1408FDC00000000000AE0BD3;
    rom[174] = 120'h0AE041D8EC33700000000AF0B63;
    rom[175] = 120'h0AF1408F6400000000000B00B33;
    rom[176] = 120'h0B01408F4400000000000B10B23;
    rom[177] = 120'h0B1300000000000000000000001;
    rom[178] = 120'h0B2300000000000000000000001;
    rom[179] = 120'h0B31408F6C00000000000B40B53;
    rom[180] = 120'h0B4300000000000000000000000;
    rom[181] = 120'h0B5300000000000000000000000;
    rom[182] = 120'h0B61408F6400000000000B70BA3;
    rom[183] = 120'h0B7A43B34813B00000000B80B93;
    rom[184] = 120'h0B8300000000000000000000001;
    rom[185] = 120'h0B9300000000000000000000000;
    rom[186] = 120'h0BAA43E1E29A000000000BB0BC3;
    rom[187] = 120'h0BB300000000000000000000000;
    rom[188] = 120'h0BC300000000000000000000001;
    rom[189] = 120'h0BD041D8EC33700000000BE0C53;
    rom[190] = 120'h0BE14094AA00000000000BF0C23;
    rom[191] = 120'h0BFA3FE00000000000000C00C13;
    rom[192] = 120'h0C0300000000000000000000000;
    rom[193] = 120'h0C1300000000000000000000001;
    rom[194] = 120'h0C21409DC200000000000C30C43;
    rom[195] = 120'h0C3300000000000000000000001;
    rom[196] = 120'h0C4300000000000000000000001;
    rom[197] = 120'h0C514094AC00000000000C60C93;
    rom[198] = 120'h0C6140930200000000000C70C83;
    rom[199] = 120'h0C7300000000000000000000001;
    rom[200] = 120'h0C8300000000000000000000001;
    rom[201] = 120'h0C91409DC200000000000CA0CB3;
    rom[202] = 120'h0CA300000000000000000000001;
    rom[203] = 120'h0CB300000000000000000000001;
    rom[204] = 120'h0CC041D8EC33B00000000CD0F03;
    rom[205] = 120'h0CDA42D00000200000000CE0E93;
    rom[206] = 120'h0CE1406BA000000000000CF0D63;
    rom[207] = 120'h0CFA419C0082100000000D00D53;
    rom[208] = 120'h0D0A40C00800000000000D10D23;
    rom[209] = 120'h0D1300000000000000000000001;
    rom[210] = 120'h0D2A418C0104200000000D30D43;
    rom[211] = 120'h0D3300000000000000000000000;
    rom[212] = 120'h0D4300000000000000000000001;
    rom[213] = 120'h0D5300000000000000000000000;
    rom[214] = 120'h0D61408CCC00000000000D70E43;
    rom[215] = 120'h0D714075F800000000000D80DF3;
    rom[216] = 120'h0D81406EA000000000000D90DA3;
    rom[217] = 120'h0D9300000000000000000000000;
    rom[218] = 120'h0DA14070C800000000000DB0DC3;
    rom[219] = 120'h0DB300000000000000000000001;
    rom[220] = 120'h0DC14073C000000000000DD0DE3;
    rom[221] = 120'h0DD300000000000000000000000;
    rom[222] = 120'h0DE300000000000000000000001;
    rom[223] = 120'h0DF1408A4800000000000E00E13;
    rom[224] = 120'h0E0300000000000000000000000;
    rom[225] = 120'h0E1A4201C199158000000E20E33;
    rom[226] = 120'h0E2300000000000000000000000;
    rom[227] = 120'h0E3300000000000000000000001;
    rom[228] = 120'h0E4A41E00000270000000E50E63;
    rom[229] = 120'h0E5300000000000000000000000;
    rom[230] = 120'h0E6A425C480B800000000E70E83;
    rom[231] = 120'h0E7300000000000000000000001;
    rom[232] = 120'h0E8300000000000000000000000;
    rom[233] = 120'h0E91407F3000000000000EA0EB3;
    rom[234] = 120'h0EA300000000000000000000000;
    rom[235] = 120'h0EBA43AA0919500000000EC0ED3;
    rom[236] = 120'h0EC300000000000000000000000;
    rom[237] = 120'h0EDA43AA7215800000000EE0EF3;
    rom[238] = 120'h0EE300000000000000000000001;
    rom[239] = 120'h0EF300000000000000000000000;
    rom[240] = 120'h0F01408EE800000000000F10F23;
    rom[241] = 120'h0F1300000000000000000000000;
    rom[242] = 120'h0F21408F5800000000000F30FC3;
    rom[243] = 120'h0F3041D8EC33D00000000F40F73;
    rom[244] = 120'h0F4A43BBF184C00000000F50F63;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
