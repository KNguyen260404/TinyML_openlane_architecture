module tree_rom_18 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000140681000000000000010023;
    rom[1] = 120'h001300000000000000000000001;
    rom[2] = 120'h002041D8EC33900000000030B43;
    rom[3] = 120'h003041D8EC33500000000040573;
    rom[4] = 120'h0041407F5800000000000050363;
    rom[5] = 120'h00514077C8000000000000601F3;
    rom[6] = 120'h006140689000000000000070103;
    rom[7] = 120'h0071406830000000000000800F3;
    rom[8] = 120'h008A4203FB67E000000000900C3;
    rom[9] = 120'h009A403700000000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00CA43D277D43000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00F300000000000000000000001;
    rom[16] = 120'h0101406F3000000000000110183;
    rom[17] = 120'h011140693000000000000120153;
    rom[18] = 120'h012A43CAD36C200000000130143;
    rom[19] = 120'h013300000000000000000000000;
    rom[20] = 120'h014300000000000000000000001;
    rom[21] = 120'h0151406E1000000000000160173;
    rom[22] = 120'h016300000000000000000000001;
    rom[23] = 120'h017300000000000000000000000;
    rom[24] = 120'h018A40B3EB800000000001901C3;
    rom[25] = 120'h019A40AF37000000000001A01B3;
    rom[26] = 120'h01A300000000000000000000001;
    rom[27] = 120'h01B300000000000000000000000;
    rom[28] = 120'h01CA43D1C0F3A000000001D01E3;
    rom[29] = 120'h01D300000000000000000000001;
    rom[30] = 120'h01E300000000000000000000001;
    rom[31] = 120'h01FA43EA3BB63000000002002F3;
    rom[32] = 120'h020A436FE816D00000000210283;
    rom[33] = 120'h021A43230018100000000220253;
    rom[34] = 120'h022A3FF80000000000000230243;
    rom[35] = 120'h023300000000000000000000000;
    rom[36] = 120'h024300000000000000000000000;
    rom[37] = 120'h0251407E8800000000000260273;
    rom[38] = 120'h026300000000000000000000001;
    rom[39] = 120'h027300000000000000000000001;
    rom[40] = 120'h0281407908000000000002902C3;
    rom[41] = 120'h029A439406C07000000002A02B3;
    rom[42] = 120'h02A300000000000000000000000;
    rom[43] = 120'h02B300000000000000000000001;
    rom[44] = 120'h02CA43D4734A1000000002D02E3;
    rom[45] = 120'h02D300000000000000000000000;
    rom[46] = 120'h02E300000000000000000000000;
    rom[47] = 120'h02F140799800000000000300353;
    rom[48] = 120'h030A43EB0586600000000310343;
    rom[49] = 120'h031A43EAD51B400000000320333;
    rom[50] = 120'h032300000000000000000000001;
    rom[51] = 120'h033300000000000000000000000;
    rom[52] = 120'h034300000000000000000000001;
    rom[53] = 120'h035300000000000000000000001;
    rom[54] = 120'h0361408FDC00000000000370463;
    rom[55] = 120'h037140861400000000000380393;
    rom[56] = 120'h038300000000000000000000001;
    rom[57] = 120'h039A3FE000000000000003A03F3;
    rom[58] = 120'h03A14088D8000000000003B03C3;
    rom[59] = 120'h03B300000000000000000000001;
    rom[60] = 120'h03C1408C58000000000003D03E3;
    rom[61] = 120'h03D300000000000000000000000;
    rom[62] = 120'h03E300000000000000000000000;
    rom[63] = 120'h03FA43A45D55300000000400433;
    rom[64] = 120'h040140861C00000000000410423;
    rom[65] = 120'h041300000000000000000000000;
    rom[66] = 120'h042300000000000000000000001;
    rom[67] = 120'h043A43E00172800000000440453;
    rom[68] = 120'h044300000000000000000000001;
    rom[69] = 120'h045300000000000000000000001;
    rom[70] = 120'h046A3FE000000000000004704E3;
    rom[71] = 120'h04714092C000000000000480493;
    rom[72] = 120'h048300000000000000000000001;
    rom[73] = 120'h0491409D06000000000004A04D3;
    rom[74] = 120'h04A140950C000000000004B04C3;
    rom[75] = 120'h04B300000000000000000000000;
    rom[76] = 120'h04C300000000000000000000001;
    rom[77] = 120'h04D300000000000000000000000;
    rom[78] = 120'h04EA43D1CCAD0000000004F0563;
    rom[79] = 120'h04F14094AA00000000000500533;
    rom[80] = 120'h050140930200000000000510523;
    rom[81] = 120'h051300000000000000000000001;
    rom[82] = 120'h052300000000000000000000001;
    rom[83] = 120'h0531409DC200000000000540553;
    rom[84] = 120'h054300000000000000000000001;
    rom[85] = 120'h055300000000000000000000001;
    rom[86] = 120'h056300000000000000000000001;
    rom[87] = 120'h057A43D3FFD9800000000580913;
    rom[88] = 120'h0581407E5800000000000590783;
    rom[89] = 120'h05914077C8000000000005A0693;
    rom[90] = 120'h05A041D8EC337000000005B0623;
    rom[91] = 120'h05BA40ADAD000000000005C05F3;
    rom[92] = 120'h05C14068C0000000000005D05E3;
    rom[93] = 120'h05D300000000000000000000000;
    rom[94] = 120'h05E300000000000000000000001;
    rom[95] = 120'h05F1406F3000000000000600613;
    rom[96] = 120'h060300000000000000000000000;
    rom[97] = 120'h061300000000000000000000001;
    rom[98] = 120'h06214068B000000000000630663;
    rom[99] = 120'h063140683000000000000640653;
    rom[100] = 120'h064300000000000000000000000;
    rom[101] = 120'h065300000000000000000000000;
    rom[102] = 120'h0661406E1000000000000670683;
    rom[103] = 120'h067300000000000000000000001;
    rom[104] = 120'h068300000000000000000000000;
    rom[105] = 120'h0691407E08000000000006A0713;
    rom[106] = 120'h06AA41EFC64F2000000006B06E3;
    rom[107] = 120'h06BA3FE000000000000006C06D3;
    rom[108] = 120'h06C300000000000000000000000;
    rom[109] = 120'h06D300000000000000000000001;
    rom[110] = 120'h06EA43B039E9A000000006F0703;
    rom[111] = 120'h06F300000000000000000000000;
    rom[112] = 120'h070300000000000000000000000;
    rom[113] = 120'h071041D8EC33700000000720753;
    rom[114] = 120'h072A41211396000000000730743;
    rom[115] = 120'h073300000000000000000000001;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h0751407E4800000000000760773;
    rom[118] = 120'h076300000000000000000000000;
    rom[119] = 120'h077300000000000000000000000;
    rom[120] = 120'h078041D8EC33700000000790883;
    rom[121] = 120'h079A3FE000000000000007A0813;
    rom[122] = 120'h07A14091AA000000000007B07E3;
    rom[123] = 120'h07B1408930000000000007C07D3;
    rom[124] = 120'h07C300000000000000000000000;
    rom[125] = 120'h07D300000000000000000000000;
    rom[126] = 120'h07E14093B4000000000007F0803;
    rom[127] = 120'h07F300000000000000000000001;
    rom[128] = 120'h080300000000000000000000000;
    rom[129] = 120'h0811408FDC00000000000820853;
    rom[130] = 120'h082A43240018100000000830843;
    rom[131] = 120'h083300000000000000000000001;
    rom[132] = 120'h084300000000000000000000001;
    rom[133] = 120'h08514094AA00000000000860873;
    rom[134] = 120'h086300000000000000000000001;
    rom[135] = 120'h087300000000000000000000001;
    rom[136] = 120'h088A3FE000000000000008908A3;
    rom[137] = 120'h089300000000000000000000000;
    rom[138] = 120'h08AA43CFF89B1000000008B08E3;
    rom[139] = 120'h08BA43AA0F0EA000000008C08D3;
    rom[140] = 120'h08C300000000000000000000001;
    rom[141] = 120'h08D300000000000000000000001;
    rom[142] = 120'h08EA43D3EE44C000000008F0903;
    rom[143] = 120'h08F300000000000000000000000;
    rom[144] = 120'h090300000000000000000000000;
    rom[145] = 120'h091041D8EC33700000000920A33;
    rom[146] = 120'h0921407F18000000000009309E3;
    rom[147] = 120'h093A43DFFC0A000000000940993;
    rom[148] = 120'h094A43D5F6CA500000000950983;
    rom[149] = 120'h095140796800000000000960973;
    rom[150] = 120'h096300000000000000000000001;
    rom[151] = 120'h097300000000000000000000001;
    rom[152] = 120'h098300000000000000000000001;
    rom[153] = 120'h0991407988000000000009A09B3;
    rom[154] = 120'h09A300000000000000000000001;
    rom[155] = 120'h09BA43EA0CFD5000000009C09D3;
    rom[156] = 120'h09C300000000000000000000000;
    rom[157] = 120'h09D300000000000000000000001;
    rom[158] = 120'h09EA43E000904000000009F0A23;
    rom[159] = 120'h09FA43DFFE83C00000000A00A13;
    rom[160] = 120'h0A0300000000000000000000001;
    rom[161] = 120'h0A1300000000000000000000000;
    rom[162] = 120'h0A2300000000000000000000001;
    rom[163] = 120'h0A31407F1800000000000A40AD3;
    rom[164] = 120'h0A4140798800000000000A50A63;
    rom[165] = 120'h0A5300000000000000000000001;
    rom[166] = 120'h0A614079E000000000000A70AA3;
    rom[167] = 120'h0A7A43EAC097800000000A80A93;
    rom[168] = 120'h0A8300000000000000000000000;
    rom[169] = 120'h0A9300000000000000000000001;
    rom[170] = 120'h0AAA43E66DE6500000000AB0AC3;
    rom[171] = 120'h0AB300000000000000000000000;
    rom[172] = 120'h0AC300000000000000000000001;
    rom[173] = 120'h0ADA43E00351200000000AE0B33;
    rom[174] = 120'h0AE1408FB000000000000AF0B23;
    rom[175] = 120'h0AF1408F6400000000000B00B13;
    rom[176] = 120'h0B0300000000000000000000001;
    rom[177] = 120'h0B1300000000000000000000000;
    rom[178] = 120'h0B2300000000000000000000001;
    rom[179] = 120'h0B3300000000000000000000001;
    rom[180] = 120'h0B4A42D00000100000000B50D63;
    rom[181] = 120'h0B5041D8EC33B00000000B60CB3;
    rom[182] = 120'h0B6A40330000000000000B70B83;
    rom[183] = 120'h0B7300000000000000000000000;
    rom[184] = 120'h0B81406BA000000000000B90C03;
    rom[185] = 120'h0B9A419C0082100000000BA0BF3;
    rom[186] = 120'h0BAA40C00800000000000BB0BC3;
    rom[187] = 120'h0BB300000000000000000000001;
    rom[188] = 120'h0BCA418C0104200000000BD0BE3;
    rom[189] = 120'h0BD300000000000000000000000;
    rom[190] = 120'h0BE300000000000000000000001;
    rom[191] = 120'h0BF300000000000000000000000;
    rom[192] = 120'h0C0A42CF8084A00000000C10C83;
    rom[193] = 120'h0C11408CCC00000000000C20C53;
    rom[194] = 120'h0C21408A4800000000000C30C43;
    rom[195] = 120'h0C3300000000000000000000000;
    rom[196] = 120'h0C4300000000000000000000000;
    rom[197] = 120'h0C5A425C480B800000000C60C73;
    rom[198] = 120'h0C6300000000000000000000001;
    rom[199] = 120'h0C7300000000000000000000000;
    rom[200] = 120'h0C814090D400000000000C90CA3;
    rom[201] = 120'h0C9300000000000000000000001;
    rom[202] = 120'h0CA300000000000000000000000;
    rom[203] = 120'h0CB041D8EC33F00000000CC0D53;
    rom[204] = 120'h0CC041D8EC33D00000000CD0CE3;
    rom[205] = 120'h0CD300000000000000000000000;
    rom[206] = 120'h0CEA421C0000000000000CF0D03;
    rom[207] = 120'h0CF300000000000000000000000;
    rom[208] = 120'h0D01408B8800000000000D10D23;
    rom[209] = 120'h0D1300000000000000000000000;
    rom[210] = 120'h0D2140917400000000000D30D43;
    rom[211] = 120'h0D3300000000000000000000000;
    rom[212] = 120'h0D4300000000000000000000000;
    rom[213] = 120'h0D5300000000000000000000000;
    rom[214] = 120'h0D6041D8EC33D00000000D70E23;
    rom[215] = 120'h0D7A43AA0919500000000D80D93;
    rom[216] = 120'h0D8300000000000000000000000;
    rom[217] = 120'h0D91407F3000000000000DA0DB3;
    rom[218] = 120'h0DA300000000000000000000000;
    rom[219] = 120'h0DBA43AA3105A00000000DC0DD3;
    rom[220] = 120'h0DC300000000000000000000001;
    rom[221] = 120'h0DD1408F5800000000000DE0E13;
    rom[222] = 120'h0DEA43BF4C03D00000000DF0E03;
    rom[223] = 120'h0DF300000000000000000000000;
    rom[224] = 120'h0E0300000000000000000000000;
    rom[225] = 120'h0E1300000000000000000000000;
    rom[226] = 120'h0E2300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 227; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
