module tree_rom_0 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    /* verilator lint_off UNUSEDSIGNAL */
    input wire [ADDR_WIDTH-1:0] addr,
    /* verilator lint_on UNUSEDSIGNAL */
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000041D8EC33900000000010B23;
    rom[1] = 120'h001140681000000000000020033;
    rom[2] = 120'h002300000000000000000000001;
    rom[3] = 120'h003A43D3FFCBB00000000040793;
    rom[4] = 120'h004A4360009A7000000000503E3;
    rom[5] = 120'h005A432318AC300000000060253;
    rom[6] = 120'h006041D8EC33500000000070163;
    rom[7] = 120'h007A417007166000000000800F3;
    rom[8] = 120'h0081406890000000000000900C3;
    rom[9] = 120'h0091406830000000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00CA3FE000000000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00FA43188B8B900000000100133;
    rom[16] = 120'h0101408A5400000000000110123;
    rom[17] = 120'h011300000000000000000000000;
    rom[18] = 120'h012300000000000000000000001;
    rom[19] = 120'h013A431D9A8AC00000000140153;
    rom[20] = 120'h014300000000000000000000000;
    rom[21] = 120'h015300000000000000000000000;
    rom[22] = 120'h0161408A54000000000001701E3;
    rom[23] = 120'h0171406E10000000000001801B3;
    rom[24] = 120'h018041D8EC337000000001901A3;
    rom[25] = 120'h019300000000000000000000001;
    rom[26] = 120'h01A300000000000000000000001;
    rom[27] = 120'h01BA400400000000000001C01D3;
    rom[28] = 120'h01C300000000000000000000000;
    rom[29] = 120'h01D300000000000000000000000;
    rom[30] = 120'h01EA3FE000000000000001F0223;
    rom[31] = 120'h01F041D8EC33700000000200213;
    rom[32] = 120'h020300000000000000000000000;
    rom[33] = 120'h021300000000000000000000000;
    rom[34] = 120'h022041D8EC33700000000230243;
    rom[35] = 120'h023300000000000000000000001;
    rom[36] = 120'h024300000000000000000000001;
    rom[37] = 120'h02514068E0000000000002602F3;
    rom[38] = 120'h026140683000000000000270283;
    rom[39] = 120'h027300000000000000000000000;
    rom[40] = 120'h028A434F1C26C000000002902C3;
    rom[41] = 120'h0291406890000000000002A02B3;
    rom[42] = 120'h02A300000000000000000000001;
    rom[43] = 120'h02B300000000000000000000000;
    rom[44] = 120'h02C1406890000000000002D02E3;
    rom[45] = 120'h02D300000000000000000000001;
    rom[46] = 120'h02E300000000000000000000000;
    rom[47] = 120'h02F041D8EC33700000000300373;
    rom[48] = 120'h030041D8EC33500000000310343;
    rom[49] = 120'h031140694000000000000320333;
    rom[50] = 120'h032300000000000000000000000;
    rom[51] = 120'h033300000000000000000000001;
    rom[52] = 120'h034A43240018100000000350363;
    rom[53] = 120'h035300000000000000000000001;
    rom[54] = 120'h036300000000000000000000001;
    rom[55] = 120'h037A4329D6A57000000003803B3;
    rom[56] = 120'h038A432585E50000000003903A3;
    rom[57] = 120'h039300000000000000000000001;
    rom[58] = 120'h03A300000000000000000000001;
    rom[59] = 120'h03BA4354B39CA000000003C03D3;
    rom[60] = 120'h03C300000000000000000000001;
    rom[61] = 120'h03D300000000000000000000001;
    rom[62] = 120'h03E041D8EC337000000003F05E3;
    rom[63] = 120'h03FA43A0B44F6000000004004F3;
    rom[64] = 120'h040041D8EC33500000000410483;
    rom[65] = 120'h041A436FE5EA600000000420453;
    rom[66] = 120'h042A436087DC400000000430443;
    rom[67] = 120'h043300000000000000000000000;
    rom[68] = 120'h044300000000000000000000001;
    rom[69] = 120'h045A4397F2DF000000000460473;
    rom[70] = 120'h046300000000000000000000000;
    rom[71] = 120'h047300000000000000000000000;
    rom[72] = 120'h0481407F70000000000004904C3;
    rom[73] = 120'h049A437001969000000004A04B3;
    rom[74] = 120'h04A300000000000000000000000;
    rom[75] = 120'h04B300000000000000000000000;
    rom[76] = 120'h04C14093C6000000000004D04E3;
    rom[77] = 120'h04D300000000000000000000001;
    rom[78] = 120'h04E300000000000000000000001;
    rom[79] = 120'h04FA43AC1BA2400000000500573;
    rom[80] = 120'h0501408F3000000000000510543;
    rom[81] = 120'h051A43A1182AA00000000520533;
    rom[82] = 120'h052300000000000000000000000;
    rom[83] = 120'h053300000000000000000000001;
    rom[84] = 120'h054041D8EC33500000000550563;
    rom[85] = 120'h055300000000000000000000001;
    rom[86] = 120'h056300000000000000000000001;
    rom[87] = 120'h0571407E98000000000005805B3;
    rom[88] = 120'h05814068B0000000000005905A3;
    rom[89] = 120'h059300000000000000000000000;
    rom[90] = 120'h05A300000000000000000000000;
    rom[91] = 120'h05BA43AE1E002000000005C05D3;
    rom[92] = 120'h05C300000000000000000000000;
    rom[93] = 120'h05D300000000000000000000001;
    rom[94] = 120'h05EA43A146635000000005F06A3;
    rom[95] = 120'h05FA437000DAE80000000600653;
    rom[96] = 120'h060A436005FE300000000610623;
    rom[97] = 120'h061300000000000000000000000;
    rom[98] = 120'h062A43607028400000000630643;
    rom[99] = 120'h063300000000000000000000001;
    rom[100] = 120'h064300000000000000000000000;
    rom[101] = 120'h06514094BC00000000000660693;
    rom[102] = 120'h066A4399A24B800000000670683;
    rom[103] = 120'h067300000000000000000000000;
    rom[104] = 120'h068300000000000000000000000;
    rom[105] = 120'h069300000000000000000000001;
    rom[106] = 120'h06A1407E98000000000006B0723;
    rom[107] = 120'h06B1407970000000000006C06F3;
    rom[108] = 120'h06CA43C21300C000000006D06E3;
    rom[109] = 120'h06D300000000000000000000000;
    rom[110] = 120'h06E300000000000000000000000;
    rom[111] = 120'h06F1407E1800000000000700713;
    rom[112] = 120'h070300000000000000000000000;
    rom[113] = 120'h071300000000000000000000000;
    rom[114] = 120'h072140930000000000000730763;
    rom[115] = 120'h0731408F3400000000000740753;
    rom[116] = 120'h074300000000000000000000001;
    rom[117] = 120'h075300000000000000000000001;
    rom[118] = 120'h07614094B200000000000770783;
    rom[119] = 120'h077300000000000000000000000;
    rom[120] = 120'h078300000000000000000000001;
    rom[121] = 120'h079041D8EC337000000007A09F3;
    rom[122] = 120'h07A1407F18000000000007B0943;
    rom[123] = 120'h07B041D8EC335000000007C08B3;
    rom[124] = 120'h07C1407988000000000007D0843;
    rom[125] = 120'h07D1406F30000000000007E0813;
    rom[126] = 120'h07E1406F10000000000007F0803;
    rom[127] = 120'h07F300000000000000000000001;
    rom[128] = 120'h080300000000000000000000000;
    rom[129] = 120'h081A43D5B884900000000820833;
    rom[130] = 120'h082300000000000000000000001;
    rom[131] = 120'h083300000000000000000000001;
    rom[132] = 120'h084A43EA3BB6300000000850883;
    rom[133] = 120'h08514079D800000000000860873;
    rom[134] = 120'h086300000000000000000000000;
    rom[135] = 120'h087300000000000000000000001;
    rom[136] = 120'h088A43EB0072B000000008908A3;
    rom[137] = 120'h089300000000000000000000001;
    rom[138] = 120'h08A300000000000000000000001;
    rom[139] = 120'h08B1407988000000000008C08D3;
    rom[140] = 120'h08C300000000000000000000001;
    rom[141] = 120'h08D14079D8000000000008E0913;
    rom[142] = 120'h08E1407998000000000008F0903;
    rom[143] = 120'h08F300000000000000000000000;
    rom[144] = 120'h090300000000000000000000000;
    rom[145] = 120'h0911407F0800000000000920933;
    rom[146] = 120'h092300000000000000000000001;
    rom[147] = 120'h093300000000000000000000000;
    rom[148] = 120'h094A43E000904000000009509E3;
    rom[149] = 120'h0951408F6C000000000009609D3;
    rom[150] = 120'h096041D8EC335000000009709A3;
    rom[151] = 120'h0971408F6400000000000980993;
    rom[152] = 120'h098300000000000000000000001;
    rom[153] = 120'h099300000000000000000000000;
    rom[154] = 120'h09AA43DFFE83C000000009B09C3;
    rom[155] = 120'h09B300000000000000000000001;
    rom[156] = 120'h09C300000000000000000000000;
    rom[157] = 120'h09D300000000000000000000001;
    rom[158] = 120'h09E300000000000000000000001;
    rom[159] = 120'h09FA43EA03DFA00000000A00B13;
    rom[160] = 120'h0A01407F1800000000000A10AA3;
    rom[161] = 120'h0A1140798000000000000A20A33;
    rom[162] = 120'h0A2300000000000000000000001;
    rom[163] = 120'h0A3A43DFDE11200000000A40A73;
    rom[164] = 120'h0A4140799800000000000A50A63;
    rom[165] = 120'h0A5300000000000000000000000;
    rom[166] = 120'h0A6300000000000000000000001;
    rom[167] = 120'h0A714079D800000000000A80A93;
    rom[168] = 120'h0A8300000000000000000000000;
    rom[169] = 120'h0A9300000000000000000000000;
    rom[170] = 120'h0AAA43E0011B900000000AB0B03;
    rom[171] = 120'h0AB1408FAC00000000000AC0AF3;
    rom[172] = 120'h0ACA43DFFD1AF00000000AD0AE3;
    rom[173] = 120'h0AD300000000000000000000001;
    rom[174] = 120'h0AE300000000000000000000000;
    rom[175] = 120'h0AF300000000000000000000001;
    rom[176] = 120'h0B0300000000000000000000001;
    rom[177] = 120'h0B1300000000000000000000001;
    rom[178] = 120'h0B21408EE800000000000B30D63;
    rom[179] = 120'h0B31406BA000000000000B40BD3;
    rom[180] = 120'h0B4041D8EC33B00000000B50BC3;
    rom[181] = 120'h0B5A419C0082100000000B60BB3;
    rom[182] = 120'h0B6A40C00800000000000B70B83;
    rom[183] = 120'h0B7300000000000000000000001;
    rom[184] = 120'h0B8A418C0104200000000B90BA3;
    rom[185] = 120'h0B9300000000000000000000000;
    rom[186] = 120'h0BA300000000000000000000001;
    rom[187] = 120'h0BB300000000000000000000000;
    rom[188] = 120'h0BC300000000000000000000000;
    rom[189] = 120'h0BDA42D00000100000000BE0CD3;
    rom[190] = 120'h0BE14075F800000000000BF0C83;
    rom[191] = 120'h0BF1406EA000000000000C00C13;
    rom[192] = 120'h0C0300000000000000000000000;
    rom[193] = 120'h0C1041D8EC33B00000000C20C73;
    rom[194] = 120'h0C2A41201209000000000C30C43;
    rom[195] = 120'h0C3300000000000000000000000;
    rom[196] = 120'h0C4A42C0002ECF8000000C50C63;
    rom[197] = 120'h0C5300000000000000000000001;
    rom[198] = 120'h0C6300000000000000000000001;
    rom[199] = 120'h0C7300000000000000000000000;
    rom[200] = 120'h0C81408A4800000000000C90CA3;
    rom[201] = 120'h0C9300000000000000000000000;
    rom[202] = 120'h0CAA4201C3DD17C000000CB0CC3;
    rom[203] = 120'h0CB300000000000000000000000;
    rom[204] = 120'h0CC300000000000000000000001;
    rom[205] = 120'h0CD1407F3000000000000CE0CF3;
    rom[206] = 120'h0CE300000000000000000000000;
    rom[207] = 120'h0CF041D8EC33B00000000D00D53;
    rom[208] = 120'h0D0A43A47300000000000D10D23;
    rom[209] = 120'h0D1300000000000000000000000;
    rom[210] = 120'h0D2A43AB1B00000000000D30D43;
    rom[211] = 120'h0D3300000000000000000000001;
    rom[212] = 120'h0D4300000000000000000000000;
    rom[213] = 120'h0D5300000000000000000000000;
    rom[214] = 120'h0D6A425D680B800000000D70DA3;
    rom[215] = 120'h0D7A41E00000270000000D80D93;
    rom[216] = 120'h0D8300000000000000000000000;
    rom[217] = 120'h0D9300000000000000000000001;
    rom[218] = 120'h0DA1408F5800000000000DB0DE3;
    rom[219] = 120'h0DBA43BBF184C00000000DC0DD3;
    rom[220] = 120'h0DC300000000000000000000000;
    rom[221] = 120'h0DD300000000000000000000001;
    rom[222] = 120'h0DE300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 223; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule

