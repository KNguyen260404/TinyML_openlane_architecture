module tree_rom_13 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000A43C2154C500000000010C23;
    rom[1] = 120'h001041D8EC33900000000020973;
    rom[2] = 120'h0021408E8C00000000000030623;
    rom[3] = 120'h003041D8EC335000000000402F3;
    rom[4] = 120'h004140689000000000000050163;
    rom[5] = 120'h005A436E8F469000000000600F3;
    rom[6] = 120'h006140681000000000000070083;
    rom[7] = 120'h007300000000000000000000001;
    rom[8] = 120'h008A4203FB67E000000000900C3;
    rom[9] = 120'h0091406830000000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00C1406830000000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00F140681000000000000100113;
    rom[16] = 120'h010300000000000000000000001;
    rom[17] = 120'h011140683000000000000120153;
    rom[18] = 120'h012A43750577000000000130143;
    rom[19] = 120'h013300000000000000000000000;
    rom[20] = 120'h014300000000000000000000000;
    rom[21] = 120'h015300000000000000000000001;
    rom[22] = 120'h016A3FE00000000000000170203;
    rom[23] = 120'h0171408C58000000000001801F3;
    rom[24] = 120'h0181408014000000000001901C3;
    rom[25] = 120'h0191407260000000000001A01B3;
    rom[26] = 120'h01A300000000000000000000000;
    rom[27] = 120'h01B300000000000000000000000;
    rom[28] = 120'h01C14088D8000000000001D01E3;
    rom[29] = 120'h01D300000000000000000000001;
    rom[30] = 120'h01E300000000000000000000000;
    rom[31] = 120'h01F300000000000000000000001;
    rom[32] = 120'h0201407E5800000000000210283;
    rom[33] = 120'h021140693000000000000220253;
    rom[34] = 120'h022140691000000000000230243;
    rom[35] = 120'h023300000000000000000000000;
    rom[36] = 120'h024300000000000000000000000;
    rom[37] = 120'h025A41EF885EE00000000260273;
    rom[38] = 120'h026300000000000000000000000;
    rom[39] = 120'h027300000000000000000000000;
    rom[40] = 120'h028A43700144C000000002902C3;
    rom[41] = 120'h029A416FBF5BF000000002A02B3;
    rom[42] = 120'h02A300000000000000000000001;
    rom[43] = 120'h02B300000000000000000000001;
    rom[44] = 120'h02C1407F58000000000002D02E3;
    rom[45] = 120'h02D300000000000000000000000;
    rom[46] = 120'h02E300000000000000000000001;
    rom[47] = 120'h02FA43AF4D385000000003004B3;
    rom[48] = 120'h030A43A13109000000000310403;
    rom[49] = 120'h031A4360009A700000000320393;
    rom[50] = 120'h032A432257EA200000000330363;
    rom[51] = 120'h033A41703921200000000340353;
    rom[52] = 120'h034300000000000000000000001;
    rom[53] = 120'h035300000000000000000000000;
    rom[54] = 120'h036041D8EC33700000000370383;
    rom[55] = 120'h037300000000000000000000001;
    rom[56] = 120'h038300000000000000000000001;
    rom[57] = 120'h039041D8EC337000000003A03D3;
    rom[58] = 120'h03AA4374AAB6F000000003B03C3;
    rom[59] = 120'h03B300000000000000000000000;
    rom[60] = 120'h03C300000000000000000000000;
    rom[61] = 120'h03D14066C0000000000003E03F3;
    rom[62] = 120'h03E300000000000000000000001;
    rom[63] = 120'h03F300000000000000000000000;
    rom[64] = 120'h040041D8EC33700000000410463;
    rom[65] = 120'h041A43ADE61B300000000420433;
    rom[66] = 120'h042300000000000000000000001;
    rom[67] = 120'h043A43AE1E00200000000440453;
    rom[68] = 120'h044300000000000000000000000;
    rom[69] = 120'h045300000000000000000000001;
    rom[70] = 120'h0461407EF0000000000004704A3;
    rom[71] = 120'h047A43ADBA3B400000000480493;
    rom[72] = 120'h048300000000000000000000001;
    rom[73] = 120'h049300000000000000000000000;
    rom[74] = 120'h04A300000000000000000000001;
    rom[75] = 120'h04B1407E98000000000004C0593;
    rom[76] = 120'h04CA43B0DE2CA000000004D0523;
    rom[77] = 120'h04D1406690000000000004E04F3;
    rom[78] = 120'h04E300000000000000000000001;
    rom[79] = 120'h04FA43AF84B4300000000500513;
    rom[80] = 120'h050300000000000000000000000;
    rom[81] = 120'h051300000000000000000000000;
    rom[82] = 120'h052A43B0E087500000000530563;
    rom[83] = 120'h053041D8EC33700000000540553;
    rom[84] = 120'h054300000000000000000000001;
    rom[85] = 120'h055300000000000000000000001;
    rom[86] = 120'h056A43BFF8BCB00000000570583;
    rom[87] = 120'h057300000000000000000000000;
    rom[88] = 120'h058300000000000000000000000;
    rom[89] = 120'h059A43C1FD881000000005A05F3;
    rom[90] = 120'h05AA43C17FEB9000000005B05C3;
    rom[91] = 120'h05B300000000000000000000001;
    rom[92] = 120'h05CA43C18BE5C000000005D05E3;
    rom[93] = 120'h05D300000000000000000000000;
    rom[94] = 120'h05E300000000000000000000001;
    rom[95] = 120'h05F14085FC00000000000600613;
    rom[96] = 120'h060300000000000000000000000;
    rom[97] = 120'h061300000000000000000000001;
    rom[98] = 120'h062A3FE000000000000006306E3;
    rom[99] = 120'h063140900200000000000640653;
    rom[100] = 120'h064300000000000000000000000;
    rom[101] = 120'h06514093B400000000000660673;
    rom[102] = 120'h066300000000000000000000001;
    rom[103] = 120'h0671409D5E000000000006806D3;
    rom[104] = 120'h068041D8EC337000000006906C3;
    rom[105] = 120'h069041D8EC335000000006A06B3;
    rom[106] = 120'h06A300000000000000000000000;
    rom[107] = 120'h06B300000000000000000000000;
    rom[108] = 120'h06C300000000000000000000000;
    rom[109] = 120'h06D300000000000000000000000;
    rom[110] = 120'h06EA426C2589E000000006F0823;
    rom[111] = 120'h06F041D8EC337000000007007B3;
    rom[112] = 120'h070041D8EC33500000000710763;
    rom[113] = 120'h0711408FDC00000000000720753;
    rom[114] = 120'h0721408FC400000000000730743;
    rom[115] = 120'h073300000000000000000000001;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h075300000000000000000000001;
    rom[118] = 120'h0761408FDC000000000007707A3;
    rom[119] = 120'h077A40A6E800000000000780793;
    rom[120] = 120'h078300000000000000000000000;
    rom[121] = 120'h079300000000000000000000001;
    rom[122] = 120'h07A300000000000000000000001;
    rom[123] = 120'h07BA408404000000000007C0813;
    rom[124] = 120'h07C1408FE4000000000007D0803;
    rom[125] = 120'h07D1408F9C000000000007E07F3;
    rom[126] = 120'h07E300000000000000000000001;
    rom[127] = 120'h07F300000000000000000000000;
    rom[128] = 120'h080300000000000000000000001;
    rom[129] = 120'h081300000000000000000000001;
    rom[130] = 120'h08214094AA00000000000830903;
    rom[131] = 120'h08314094A6000000000008408B3;
    rom[132] = 120'h084041D8EC33700000000850883;
    rom[133] = 120'h0851408FCC00000000000860873;
    rom[134] = 120'h086300000000000000000000000;
    rom[135] = 120'h087300000000000000000000001;
    rom[136] = 120'h088A43B33A1D7000000008908A3;
    rom[137] = 120'h089300000000000000000000000;
    rom[138] = 120'h08A300000000000000000000001;
    rom[139] = 120'h08B041D8EC337000000008C08F3;
    rom[140] = 120'h08C041D8EC335000000008D08E3;
    rom[141] = 120'h08D300000000000000000000000;
    rom[142] = 120'h08E300000000000000000000000;
    rom[143] = 120'h08F300000000000000000000000;
    rom[144] = 120'h090A42D0011EF00000000910963;
    rom[145] = 120'h091A42CFFE12900000000920953;
    rom[146] = 120'h092A42C3FCDDC00000000930943;
    rom[147] = 120'h093300000000000000000000001;
    rom[148] = 120'h094300000000000000000000001;
    rom[149] = 120'h095300000000000000000000000;
    rom[150] = 120'h096300000000000000000000001;
    rom[151] = 120'h0971408EE800000000000980B33;
    rom[152] = 120'h0981406BA000000000000990A03;
    rom[153] = 120'h099A419C00821000000009A09F3;
    rom[154] = 120'h09AA40C008000000000009B09C3;
    rom[155] = 120'h09B300000000000000000000001;
    rom[156] = 120'h09CA418C01042000000009D09E3;
    rom[157] = 120'h09D300000000000000000000000;
    rom[158] = 120'h09E300000000000000000000001;
    rom[159] = 120'h09F300000000000000000000000;
    rom[160] = 120'h0A0A42D00000100000000A10AC3;
    rom[161] = 120'h0A1041D8EC33B00000000A20AB3;
    rom[162] = 120'h0A2A42C40000000000000A30AA3;
    rom[163] = 120'h0A31408A4800000000000A40A73;
    rom[164] = 120'h0A4A41300913000000000A50A63;
    rom[165] = 120'h0A5300000000000000000000000;
    rom[166] = 120'h0A6300000000000000000000000;
    rom[167] = 120'h0A7A4201C1B515C000000A80A93;
    rom[168] = 120'h0A8300000000000000000000000;
    rom[169] = 120'h0A9300000000000000000000001;
    rom[170] = 120'h0AA300000000000000000000001;
    rom[171] = 120'h0AB300000000000000000000000;
    rom[172] = 120'h0ACA43A56708900000000AD0AE3;
    rom[173] = 120'h0AD300000000000000000000000;
    rom[174] = 120'h0AE1407EF000000000000AF0B03;
    rom[175] = 120'h0AF300000000000000000000000;
    rom[176] = 120'h0B0A43AB1B00000000000B10B23;
    rom[177] = 120'h0B1300000000000000000000001;
    rom[178] = 120'h0B2300000000000000000000000;
    rom[179] = 120'h0B3A425D680B800000000B40B93;
    rom[180] = 120'h0B41408F9000000000000B50B83;
    rom[181] = 120'h0B5A41E00000000000000B60B73;
    rom[182] = 120'h0B6300000000000000000000000;
    rom[183] = 120'h0B7300000000000000000000001;
    rom[184] = 120'h0B8300000000000000000000000;
    rom[185] = 120'h0B9041D8EC33D00000000BA0C13;
    rom[186] = 120'h0BA041D8EC33B00000000BB0BC3;
    rom[187] = 120'h0BB300000000000000000000000;
    rom[188] = 120'h0BC1408F6800000000000BD0C03;
    rom[189] = 120'h0BDA43BBF184000000000BE0BF3;
    rom[190] = 120'h0BE300000000000000000000000;
    rom[191] = 120'h0BF300000000000000000000001;
    rom[192] = 120'h0C0300000000000000000000000;
    rom[193] = 120'h0C1300000000000000000000000;
    rom[194] = 120'h0C2A43C7FFB4800000000C30C43;
    rom[195] = 120'h0C3300000000000000000000001;
    rom[196] = 120'h0C4A43D3FFE4D00000000C51063;
    rom[197] = 120'h0C51407E9800000000000C60EF3;
    rom[198] = 120'h0C6041D8EC33700000000C70E03;
    rom[199] = 120'h0C7A43D17E79E00000000C80D73;
    rom[200] = 120'h0C8A43CA02A2600000000C90D03;
    rom[201] = 120'h0C9041D8EC33500000000CA0CD3;
    rom[202] = 120'h0CAA43C83658300000000CB0CC3;
    rom[203] = 120'h0CB300000000000000000000000;
    rom[204] = 120'h0CC300000000000000000000000;
    rom[205] = 120'h0CD14068D000000000000CE0CF3;
    rom[206] = 120'h0CE300000000000000000000000;
    rom[207] = 120'h0CF300000000000000000000001;
    rom[208] = 120'h0D0041D8EC33500000000D10D43;
    rom[209] = 120'h0D114079C800000000000D20D33;
    rom[210] = 120'h0D2300000000000000000000001;
    rom[211] = 120'h0D3300000000000000000000000;
    rom[212] = 120'h0D414079C800000000000D50D63;
    rom[213] = 120'h0D5300000000000000000000001;
    rom[214] = 120'h0D6300000000000000000000000;
    rom[215] = 120'h0D7140728800000000000D80D93;
    rom[216] = 120'h0D8300000000000000000000001;
    rom[217] = 120'h0D91407E3800000000000DA0DD3;
    rom[218] = 120'h0DA041D8EC33500000000DB0DC3;
    rom[219] = 120'h0DB300000000000000000000000;
    rom[220] = 120'h0DC300000000000000000000000;
    rom[221] = 120'h0DD1407E6800000000000DE0DF3;
    rom[222] = 120'h0DE300000000000000000000000;
    rom[223] = 120'h0DF300000000000000000000000;
    rom[224] = 120'h0E014067E000000000000E10E23;
    rom[225] = 120'h0E1300000000000000000000001;
    rom[226] = 120'h0E2A43CFE25DD00000000E30E83;
    rom[227] = 120'h0E3A43CA00A9C00000000E40E73;
    rom[228] = 120'h0E4A43C9DB9D800000000E50E63;
    rom[229] = 120'h0E5300000000000000000000000;
    rom[230] = 120'h0E6300000000000000000000000;
    rom[231] = 120'h0E7300000000000000000000001;
    rom[232] = 120'h0E8A43D17F22D00000000E90EC3;
    rom[233] = 120'h0E9A43D02BDCB00000000EA0EB3;
    rom[234] = 120'h0EA300000000000000000000000;
    rom[235] = 120'h0EB300000000000000000000001;
    rom[236] = 120'h0ECA43D1CAC4300000000ED0EE3;
    rom[237] = 120'h0ED300000000000000000000000;
    rom[238] = 120'h0EE300000000000000000000000;
    rom[239] = 120'h0EFA43D007FE700000000F00F13;
    rom[240] = 120'h0F0300000000000000000000001;
    rom[241] = 120'h0F1041D8EC33700000000F20FF3;
    rom[242] = 120'h0F2A43D013C5F00000000F30F83;
    rom[243] = 120'h0F314092A400000000000F40F53;
    rom[244] = 120'h0F4300000000000000000000001;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
