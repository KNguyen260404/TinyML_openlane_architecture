module tree_rom_7 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000041D8EC33900000000010A03;
    rom[1] = 120'h001140681000000000000020033;
    rom[2] = 120'h002300000000000000000000001;
    rom[3] = 120'h003A43D3FFE4D000000000406F3;
    rom[4] = 120'h0041407E5800000000000050403;
    rom[5] = 120'h005041D8EC33500000000060213;
    rom[6] = 120'h006A40F00178000000000070143;
    rom[7] = 120'h007A406FD0000000000000800F3;
    rom[8] = 120'h00814077E8000000000000900C3;
    rom[9] = 120'h009A3FF000000000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00C1407CD8000000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00FA40D04A40000000000100133;
    rom[16] = 120'h010A40B08600000000000110123;
    rom[17] = 120'h011300000000000000000000000;
    rom[18] = 120'h012300000000000000000000000;
    rom[19] = 120'h013300000000000000000000001;
    rom[20] = 120'h0141406930000000000001501C3;
    rom[21] = 120'h015A43CA7D45B00000000160193;
    rom[22] = 120'h016140683000000000000170183;
    rom[23] = 120'h017300000000000000000000000;
    rom[24] = 120'h018300000000000000000000000;
    rom[25] = 120'h019A43CC0B3A5000000001A01B3;
    rom[26] = 120'h01A300000000000000000000001;
    rom[27] = 120'h01B300000000000000000000001;
    rom[28] = 120'h01C1406E10000000000001D01E3;
    rom[29] = 120'h01D300000000000000000000001;
    rom[30] = 120'h01E1407838000000000001F0203;
    rom[31] = 120'h01F300000000000000000000000;
    rom[32] = 120'h020300000000000000000000000;
    rom[33] = 120'h02114077C800000000000220313;
    rom[34] = 120'h02214068B0000000000002302A3;
    rom[35] = 120'h023140689000000000000240273;
    rom[36] = 120'h024041D8EC33700000000250263;
    rom[37] = 120'h025300000000000000000000000;
    rom[38] = 120'h026300000000000000000000000;
    rom[39] = 120'h027A42000205C85C00000280293;
    rom[40] = 120'h028300000000000000000000000;
    rom[41] = 120'h029300000000000000000000000;
    rom[42] = 120'h02AA40AFDC000000000002B02E3;
    rom[43] = 120'h02B041D8EC337000000002C02D3;
    rom[44] = 120'h02C300000000000000000000001;
    rom[45] = 120'h02D300000000000000000000001;
    rom[46] = 120'h02E041D8EC337000000002F0303;
    rom[47] = 120'h02F300000000000000000000000;
    rom[48] = 120'h030300000000000000000000000;
    rom[49] = 120'h031A41EF977F200000000320393;
    rom[50] = 120'h0321407CC800000000000330363;
    rom[51] = 120'h033A413ED1EF800000000340353;
    rom[52] = 120'h034300000000000000000000000;
    rom[53] = 120'h035300000000000000000000001;
    rom[54] = 120'h0361407CD800000000000370383;
    rom[55] = 120'h037300000000000000000000000;
    rom[56] = 120'h038300000000000000000000000;
    rom[57] = 120'h039A43D17F22D000000003A03D3;
    rom[58] = 120'h03A1407C78000000000003B03C3;
    rom[59] = 120'h03B300000000000000000000000;
    rom[60] = 120'h03C300000000000000000000000;
    rom[61] = 120'h03D1407970000000000003E03F3;
    rom[62] = 120'h03E300000000000000000000001;
    rom[63] = 120'h03F300000000000000000000000;
    rom[64] = 120'h040041D8EC337000000004105E3;
    rom[65] = 120'h041A3FE000000000000004204F3;
    rom[66] = 120'h0421409002000000000004304A3;
    rom[67] = 120'h04314088D800000000000440473;
    rom[68] = 120'h044041D8EC33500000000450463;
    rom[69] = 120'h045300000000000000000000000;
    rom[70] = 120'h046300000000000000000000000;
    rom[71] = 120'h0471408C5800000000000480493;
    rom[72] = 120'h048300000000000000000000000;
    rom[73] = 120'h049300000000000000000000000;
    rom[74] = 120'h04A1409D5E000000000004B04E3;
    rom[75] = 120'h04B1409436000000000004C04D3;
    rom[76] = 120'h04C300000000000000000000000;
    rom[77] = 120'h04D300000000000000000000001;
    rom[78] = 120'h04E300000000000000000000000;
    rom[79] = 120'h04F041D8EC33500000000500573;
    rom[80] = 120'h0501408FDC00000000000510543;
    rom[81] = 120'h051A436FE82AC00000000520533;
    rom[82] = 120'h052300000000000000000000001;
    rom[83] = 120'h053300000000000000000000000;
    rom[84] = 120'h05414094AA00000000000550563;
    rom[85] = 120'h055300000000000000000000001;
    rom[86] = 120'h056300000000000000000000001;
    rom[87] = 120'h057A41701EE69800000005805B3;
    rom[88] = 120'h0581408FDC000000000005905A3;
    rom[89] = 120'h059300000000000000000000001;
    rom[90] = 120'h05A300000000000000000000001;
    rom[91] = 120'h05BA41A88EEB7000000005C05D3;
    rom[92] = 120'h05C300000000000000000000000;
    rom[93] = 120'h05D300000000000000000000001;
    rom[94] = 120'h05EA3FE000000000000005F0603;
    rom[95] = 120'h05F300000000000000000000000;
    rom[96] = 120'h060A43CFF89B100000000610683;
    rom[97] = 120'h061A43A94BD2300000000620653;
    rom[98] = 120'h062A436A870CA00000000630643;
    rom[99] = 120'h063300000000000000000000001;
    rom[100] = 120'h064300000000000000000000000;
    rom[101] = 120'h065A43AE2B12000000000660673;
    rom[102] = 120'h066300000000000000000000001;
    rom[103] = 120'h067300000000000000000000001;
    rom[104] = 120'h0681407FB8000000000006906C3;
    rom[105] = 120'h0691407E88000000000006A06B3;
    rom[106] = 120'h06A300000000000000000000001;
    rom[107] = 120'h06B300000000000000000000000;
    rom[108] = 120'h06CA43D01B853000000006D06E3;
    rom[109] = 120'h06D300000000000000000000000;
    rom[110] = 120'h06E300000000000000000000001;
    rom[111] = 120'h06FA43DEDBB4700000000700813;
    rom[112] = 120'h07014079D800000000000710803;
    rom[113] = 120'h07114079C8000000000007207D3;
    rom[114] = 120'h072140798800000000000730783;
    rom[115] = 120'h073A43D5BA8DF00000000740753;
    rom[116] = 120'h074300000000000000000000001;
    rom[117] = 120'h075041D8EC33500000000760773;
    rom[118] = 120'h076300000000000000000000001;
    rom[119] = 120'h077300000000000000000000001;
    rom[120] = 120'h078A43D5FF244000000007907C3;
    rom[121] = 120'h079A43D58F4EF000000007A07B3;
    rom[122] = 120'h07A300000000000000000000001;
    rom[123] = 120'h07B300000000000000000000000;
    rom[124] = 120'h07C300000000000000000000001;
    rom[125] = 120'h07DA43D576E0B000000007E07F3;
    rom[126] = 120'h07E300000000000000000000000;
    rom[127] = 120'h07F300000000000000000000001;
    rom[128] = 120'h080300000000000000000000001;
    rom[129] = 120'h081A43E00015900000000820913;
    rom[130] = 120'h082041D8EC337000000008308A3;
    rom[131] = 120'h083A43DFFF61A00000000840893;
    rom[132] = 120'h084041D8EC33500000000850883;
    rom[133] = 120'h0851406F6000000000000860873;
    rom[134] = 120'h086300000000000000000000000;
    rom[135] = 120'h087300000000000000000000001;
    rom[136] = 120'h088300000000000000000000001;
    rom[137] = 120'h089300000000000000000000000;
    rom[138] = 120'h08A140900C000000000008B0903;
    rom[139] = 120'h08B1407878000000000008C08D3;
    rom[140] = 120'h08C300000000000000000000001;
    rom[141] = 120'h08DA43DFFAB04000000008E08F3;
    rom[142] = 120'h08E300000000000000000000001;
    rom[143] = 120'h08F300000000000000000000000;
    rom[144] = 120'h090300000000000000000000001;
    rom[145] = 120'h0911407F18000000000009209F3;
    rom[146] = 120'h092041D8EC337000000009309A3;
    rom[147] = 120'h093041D8EC33500000000940973;
    rom[148] = 120'h094A43EA3790A00000000950963;
    rom[149] = 120'h095300000000000000000000000;
    rom[150] = 120'h096300000000000000000000001;
    rom[151] = 120'h097A43EA0545F00000000980993;
    rom[152] = 120'h098300000000000000000000000;
    rom[153] = 120'h099300000000000000000000001;
    rom[154] = 120'h09A1407988000000000009B09C3;
    rom[155] = 120'h09B300000000000000000000001;
    rom[156] = 120'h09C14079D8000000000009D09E3;
    rom[157] = 120'h09D300000000000000000000000;
    rom[158] = 120'h09E300000000000000000000000;
    rom[159] = 120'h09F300000000000000000000001;
    rom[160] = 120'h0A0041D8EC33B00000000A10C23;
    rom[161] = 120'h0A1A42D00000200000000A20BD3;
    rom[162] = 120'h0A2A40330000000000000A30A43;
    rom[163] = 120'h0A3300000000000000000000000;
    rom[164] = 120'h0A41406BA000000000000A50AC3;
    rom[165] = 120'h0A5A419C0082100000000A60AB3;
    rom[166] = 120'h0A6A40C00800000000000A70A83;
    rom[167] = 120'h0A7300000000000000000000001;
    rom[168] = 120'h0A8A418C0104200000000A90AA3;
    rom[169] = 120'h0A9300000000000000000000000;
    rom[170] = 120'h0AA300000000000000000000001;
    rom[171] = 120'h0AB300000000000000000000000;
    rom[172] = 120'h0AC1408CCC00000000000AD0B83;
    rom[173] = 120'h0AD140762000000000000AE0B33;
    rom[174] = 120'h0AEA42C0002ECF8000000AF0B23;
    rom[175] = 120'h0AFA41944607920000000B00B13;
    rom[176] = 120'h0B0300000000000000000000000;
    rom[177] = 120'h0B1300000000000000000000000;
    rom[178] = 120'h0B2300000000000000000000001;
    rom[179] = 120'h0B3A420D9010E00000000B40B53;
    rom[180] = 120'h0B4300000000000000000000000;
    rom[181] = 120'h0B5140890C00000000000B60B73;
    rom[182] = 120'h0B6300000000000000000000000;
    rom[183] = 120'h0B7300000000000000000000001;
    rom[184] = 120'h0B81408F9000000000000B90BC3;
    rom[185] = 120'h0B9A42651000400000000BA0BB3;
    rom[186] = 120'h0BA300000000000000000000001;
    rom[187] = 120'h0BB300000000000000000000000;
    rom[188] = 120'h0BC300000000000000000000000;
    rom[189] = 120'h0BDA43AA8E01C00000000BE0C13;
    rom[190] = 120'h0BEA43AA0919500000000BF0C03;
    rom[191] = 120'h0BF300000000000000000000000;
    rom[192] = 120'h0C0300000000000000000000001;
    rom[193] = 120'h0C1300000000000000000000000;
    rom[194] = 120'h0C2A43BBF184C00000000C30CE3;
    rom[195] = 120'h0C3041D8EC33F00000000C40CD3;
    rom[196] = 120'h0C4041D8EC33D00000000C50C63;
    rom[197] = 120'h0C5300000000000000000000000;
    rom[198] = 120'h0C6A42250000000000000C70CC3;
    rom[199] = 120'h0C71408CCC00000000000C80C93;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C9A42140000040000000CA0CB3;
    rom[202] = 120'h0CA300000000000000000000000;
    rom[203] = 120'h0CB300000000000000000000001;
    rom[204] = 120'h0CC300000000000000000000000;
    rom[205] = 120'h0CD300000000000000000000000;
    rom[206] = 120'h0CE140877800000000000CF0D03;
    rom[207] = 120'h0CF300000000000000000000000;
    rom[208] = 120'h0D0041D8EC33D00000000D10D43;
    rom[209] = 120'h0D1A43C02A4F380000000D20D33;
    rom[210] = 120'h0D2300000000000000000000001;
    rom[211] = 120'h0D3300000000000000000000000;
    rom[212] = 120'h0D4300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 213; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
