module tree_rom_10 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000041D8EC33900000000011083;
    rom[1] = 120'h001A43C2154BD00000000020B73;
    rom[2] = 120'h002041D8EC33500000000030503;
    rom[3] = 120'h003A41701FB2800000000040273;
    rom[4] = 120'h004A4136BE2B8000000000501A3;
    rom[5] = 120'h0051406890000000000000600B3;
    rom[6] = 120'h006140681000000000000070083;
    rom[7] = 120'h007300000000000000000000001;
    rom[8] = 120'h008A403700000000000000900A3;
    rom[9] = 120'h009300000000000000000000001;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00BA3FE000000000000000C0133;
    rom[12] = 120'h00C1409002000000000000D0103;
    rom[13] = 120'h00D1408C58000000000000E00F3;
    rom[14] = 120'h00E300000000000000000000000;
    rom[15] = 120'h00F300000000000000000000000;
    rom[16] = 120'h01014092C000000000000110123;
    rom[17] = 120'h011300000000000000000000001;
    rom[18] = 120'h012300000000000000000000000;
    rom[19] = 120'h0131407E1800000000000140173;
    rom[20] = 120'h014A40F00178000000000150163;
    rom[21] = 120'h015300000000000000000000001;
    rom[22] = 120'h016300000000000000000000000;
    rom[23] = 120'h0171408FDC00000000000180193;
    rom[24] = 120'h018300000000000000000000001;
    rom[25] = 120'h019300000000000000000000001;
    rom[26] = 120'h01A1408A5C000000000001B0263;
    rom[27] = 120'h01B1408A3C000000000001C0213;
    rom[28] = 120'h01C14079E0000000000001D0203;
    rom[29] = 120'h01D14079C8000000000001E01F3;
    rom[30] = 120'h01E300000000000000000000001;
    rom[31] = 120'h01F300000000000000000000000;
    rom[32] = 120'h020300000000000000000000001;
    rom[33] = 120'h0211408A4400000000000220233;
    rom[34] = 120'h022300000000000000000000000;
    rom[35] = 120'h0231408A4C00000000000240253;
    rom[36] = 120'h024300000000000000000000001;
    rom[37] = 120'h025300000000000000000000000;
    rom[38] = 120'h026300000000000000000000001;
    rom[39] = 120'h0271407E5800000000000280393;
    rom[40] = 120'h0281406810000000000002902A3;
    rom[41] = 120'h029300000000000000000000001;
    rom[42] = 120'h02AA41EF934BC000000002B0323;
    rom[43] = 120'h02B1406E10000000000002C02F3;
    rom[44] = 120'h02C1406950000000000002D02E3;
    rom[45] = 120'h02D300000000000000000000000;
    rom[46] = 120'h02E300000000000000000000001;
    rom[47] = 120'h02FA41DFCE58400000000300313;
    rom[48] = 120'h030300000000000000000000000;
    rom[49] = 120'h031300000000000000000000001;
    rom[50] = 120'h032140693000000000000330363;
    rom[51] = 120'h033A4209FAFC400000000340353;
    rom[52] = 120'h034300000000000000000000001;
    rom[53] = 120'h035300000000000000000000000;
    rom[54] = 120'h036A43B1CC90D00000000370383;
    rom[55] = 120'h037300000000000000000000000;
    rom[56] = 120'h038300000000000000000000001;
    rom[57] = 120'h0391408FCC000000000003A0473;
    rom[58] = 120'h03AA436FE82AC000000003B0423;
    rom[59] = 120'h03BA42A26B7A1000000003C03F3;
    rom[60] = 120'h03C1408A54000000000003D03E3;
    rom[61] = 120'h03D300000000000000000000000;
    rom[62] = 120'h03E300000000000000000000001;
    rom[63] = 120'h03F1408F4000000000000400413;
    rom[64] = 120'h040300000000000000000000001;
    rom[65] = 120'h041300000000000000000000000;
    rom[66] = 120'h042A43B01A13B80000000430463;
    rom[67] = 120'h043A43AE1616700000000440453;
    rom[68] = 120'h044300000000000000000000000;
    rom[69] = 120'h045300000000000000000000000;
    rom[70] = 120'h046300000000000000000000001;
    rom[71] = 120'h047A43C20FC12000000004804F3;
    rom[72] = 120'h04814093C6000000000004904C3;
    rom[73] = 120'h049A426C19A90000000004A04B3;
    rom[74] = 120'h04A300000000000000000000001;
    rom[75] = 120'h04B300000000000000000000001;
    rom[76] = 120'h04CA42D0011EF000000004D04E3;
    rom[77] = 120'h04D300000000000000000000001;
    rom[78] = 120'h04E300000000000000000000001;
    rom[79] = 120'h04F300000000000000000000000;
    rom[80] = 120'h050041D8EC337000000005108C3;
    rom[81] = 120'h051A436000A11000000005206F3;
    rom[82] = 120'h052A4323ED19000000000530623;
    rom[83] = 120'h053A42EFFD50F000000005405B3;
    rom[84] = 120'h0541408A5400000000000550583;
    rom[85] = 120'h055A41703921200000000560573;
    rom[86] = 120'h056300000000000000000000001;
    rom[87] = 120'h057300000000000000000000000;
    rom[88] = 120'h058A3FE000000000000005905A3;
    rom[89] = 120'h059300000000000000000000000;
    rom[90] = 120'h05A300000000000000000000001;
    rom[91] = 120'h05B1407F38000000000005C05F3;
    rom[92] = 120'h05CA431C60169000000005D05E3;
    rom[93] = 120'h05D300000000000000000000000;
    rom[94] = 120'h05E300000000000000000000000;
    rom[95] = 120'h05F140907A00000000000600613;
    rom[96] = 120'h060300000000000000000000001;
    rom[97] = 120'h061300000000000000000000001;
    rom[98] = 120'h06214068D0000000000006306A3;
    rom[99] = 120'h063A4340B26D000000000640673;
    rom[100] = 120'h064A433C6AAE000000000650663;
    rom[101] = 120'h065300000000000000000000001;
    rom[102] = 120'h066300000000000000000000001;
    rom[103] = 120'h067A434D0C03A00000000680693;
    rom[104] = 120'h068300000000000000000000000;
    rom[105] = 120'h069300000000000000000000000;
    rom[106] = 120'h06A1407E80000000000006B06C3;
    rom[107] = 120'h06B300000000000000000000001;
    rom[108] = 120'h06C1408FD0000000000006D06E3;
    rom[109] = 120'h06D300000000000000000000001;
    rom[110] = 120'h06E300000000000000000000001;
    rom[111] = 120'h06FA43A100689000000007007D3;
    rom[112] = 120'h0701407F7000000000000710763;
    rom[113] = 120'h071140681000000000000720733;
    rom[114] = 120'h072300000000000000000000001;
    rom[115] = 120'h0731406EF000000000000740753;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h075300000000000000000000000;
    rom[118] = 120'h0761408F8C000000000007707A3;
    rom[119] = 120'h077A439D7F95700000000780793;
    rom[120] = 120'h078300000000000000000000001;
    rom[121] = 120'h079300000000000000000000000;
    rom[122] = 120'h07AA439FCC80D000000007B07C3;
    rom[123] = 120'h07B300000000000000000000001;
    rom[124] = 120'h07C300000000000000000000000;
    rom[125] = 120'h07DA43AE0DD79000000007E0853;
    rom[126] = 120'h07EA43A514B2E000000007F0823;
    rom[127] = 120'h07FA43A11896E00000000800813;
    rom[128] = 120'h080300000000000000000000000;
    rom[129] = 120'h081300000000000000000000001;
    rom[130] = 120'h0821408F3000000000000830843;
    rom[131] = 120'h083300000000000000000000001;
    rom[132] = 120'h084300000000000000000000001;
    rom[133] = 120'h085A43B0E066D00000000860893;
    rom[134] = 120'h0861407F6000000000000870883;
    rom[135] = 120'h087300000000000000000000000;
    rom[136] = 120'h088300000000000000000000001;
    rom[137] = 120'h089A43BFFB011000000008A08B3;
    rom[138] = 120'h08A300000000000000000000001;
    rom[139] = 120'h08B300000000000000000000000;
    rom[140] = 120'h08C1407E18000000000008D0A23;
    rom[141] = 120'h08DA40F7FDD80000000008E0993;
    rom[142] = 120'h08E1407328000000000008F0943;
    rom[143] = 120'h08F1406DE000000000000900913;
    rom[144] = 120'h090300000000000000000000001;
    rom[145] = 120'h0911406E8000000000000920933;
    rom[146] = 120'h092300000000000000000000000;
    rom[147] = 120'h093300000000000000000000001;
    rom[148] = 120'h0941407CF000000000000950983;
    rom[149] = 120'h0951407CC800000000000960973;
    rom[150] = 120'h096300000000000000000000000;
    rom[151] = 120'h097300000000000000000000000;
    rom[152] = 120'h098300000000000000000000001;
    rom[153] = 120'h0991406810000000000009A09B3;
    rom[154] = 120'h09A300000000000000000000001;
    rom[155] = 120'h09BA436080074000000009C09F3;
    rom[156] = 120'h09C1407838000000000009D09E3;
    rom[157] = 120'h09D300000000000000000000000;
    rom[158] = 120'h09E300000000000000000000000;
    rom[159] = 120'h09F1407C3800000000000A00A13;
    rom[160] = 120'h0A0300000000000000000000000;
    rom[161] = 120'h0A1300000000000000000000001;
    rom[162] = 120'h0A2140861400000000000A30AC3;
    rom[163] = 120'h0A3A3FF00000000000000A40A53;
    rom[164] = 120'h0A4300000000000000000000000;
    rom[165] = 120'h0A51407E9800000000000A60A93;
    rom[166] = 120'h0A61407E8000000000000A70A83;
    rom[167] = 120'h0A7300000000000000000000001;
    rom[168] = 120'h0A8300000000000000000000001;
    rom[169] = 120'h0A91407F5800000000000AA0AB3;
    rom[170] = 120'h0AA300000000000000000000001;
    rom[171] = 120'h0AB300000000000000000000001;
    rom[172] = 120'h0AC1408E9000000000000AD0B23;
    rom[173] = 120'h0ADA439DD3FEC00000000AE0B13;
    rom[174] = 120'h0AE1408A5C00000000000AF0B03;
    rom[175] = 120'h0AF300000000000000000000000;
    rom[176] = 120'h0B0300000000000000000000000;
    rom[177] = 120'h0B1300000000000000000000001;
    rom[178] = 120'h0B2A3FF00000000000000B30B43;
    rom[179] = 120'h0B3300000000000000000000000;
    rom[180] = 120'h0B41408F8000000000000B50B63;
    rom[181] = 120'h0B5300000000000000000000001;
    rom[182] = 120'h0B6300000000000000000000001;
    rom[183] = 120'h0B7A43C7FFA6C00000000B80B93;
    rom[184] = 120'h0B8300000000000000000000001;
    rom[185] = 120'h0B9041D8EC33700000000BA0E73;
    rom[186] = 120'h0BA1407F1800000000000BB0D83;
    rom[187] = 120'h0BB140798800000000000BC0C93;
    rom[188] = 120'h0BC041D8EC33500000000BD0C23;
    rom[189] = 120'h0BD14072A800000000000BE0C13;
    rom[190] = 120'h0BEA43CA027DA00000000BF0C03;
    rom[191] = 120'h0BF300000000000000000000000;
    rom[192] = 120'h0C0300000000000000000000001;
    rom[193] = 120'h0C1300000000000000000000001;
    rom[194] = 120'h0C2A43CA14FBE00000000C30C63;
    rom[195] = 120'h0C3140676000000000000C40C53;
    rom[196] = 120'h0C4300000000000000000000001;
    rom[197] = 120'h0C5300000000000000000000000;
    rom[198] = 120'h0C6A43D1C6E0700000000C70C83;
    rom[199] = 120'h0C7300000000000000000000001;
    rom[200] = 120'h0C8300000000000000000000001;
    rom[201] = 120'h0C9A43EA3A6F100000000CA0D13;
    rom[202] = 120'h0CAA43D40221F00000000CB0CE3;
    rom[203] = 120'h0CBA43CFF997D00000000CC0CD3;
    rom[204] = 120'h0CC300000000000000000000001;
    rom[205] = 120'h0CD300000000000000000000000;
    rom[206] = 120'h0CE041D8EC33500000000CF0D03;
    rom[207] = 120'h0CF300000000000000000000000;
    rom[208] = 120'h0D0300000000000000000000000;
    rom[209] = 120'h0D1041D8EC33500000000D20D53;
    rom[210] = 120'h0D214079A000000000000D30D43;
    rom[211] = 120'h0D3300000000000000000000000;
    rom[212] = 120'h0D4300000000000000000000001;
    rom[213] = 120'h0D5A43EB03CD700000000D60D73;
    rom[214] = 120'h0D6300000000000000000000001;
    rom[215] = 120'h0D7300000000000000000000001;
    rom[216] = 120'h0D8041D8EC33500000000D90E03;
    rom[217] = 120'h0D9140945200000000000DA0DF3;
    rom[218] = 120'h0DA1408F6400000000000DB0DC3;
    rom[219] = 120'h0DB300000000000000000000001;
    rom[220] = 120'h0DC1408F6C00000000000DD0DE3;
    rom[221] = 120'h0DD300000000000000000000000;
    rom[222] = 120'h0DE300000000000000000000001;
    rom[223] = 120'h0DF300000000000000000000001;
    rom[224] = 120'h0E0A43E0009EA00000000E10E63;
    rom[225] = 120'h0E1A43DFFE83C00000000E20E53;
    rom[226] = 120'h0E2140945200000000000E30E43;
    rom[227] = 120'h0E3300000000000000000000001;
    rom[228] = 120'h0E4300000000000000000000001;
    rom[229] = 120'h0E5300000000000000000000000;
    rom[230] = 120'h0E6300000000000000000000001;
    rom[231] = 120'h0E7A43D3FFD9800000000E80F93;
    rom[232] = 120'h0E8A43CFF1FD9000000000E90F03;
    rom[233] = 120'h0E9140697000000000000EA0EF3;
    rom[234] = 120'h0EAA43CA35FF1000000000EB0EE3;
    rom[235] = 120'h0EBA43C809B3500000000EC0ED3;
    rom[236] = 120'h0EC300000000000000000000000;
    rom[237] = 120'h0ED300000000000000000000000;
    rom[238] = 120'h0EE300000000000000000000001;
    rom[239] = 120'h0EF300000000000000000000001;
    rom[240] = 120'h0F0140945C00000000000F10F83;
    rom[241] = 120'h0F1A43D1D300B00000000F20F53;
    rom[242] = 120'h0F2140729000000000000F30F43;
    rom[243] = 120'h0F3300000000000000000000001;
    rom[244] = 120'h0F4300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
