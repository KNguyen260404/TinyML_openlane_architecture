module tree_rom_14 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000140681000000000000010023;
    rom[1] = 120'h001300000000000000000000001;
    rom[2] = 120'h0021407F3800000000000030783;
    rom[3] = 120'h003041D8EC33900000000040633;
    rom[4] = 120'h00414077C8000000000000502E3;
    rom[5] = 120'h005140734800000000000060233;
    rom[6] = 120'h006A40AFDC00000000000070143;
    rom[7] = 120'h007A3FE000000000000000800F3;
    rom[8] = 120'h0081406860000000000000900C3;
    rom[9] = 120'h009041D8EC335000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000000;
    rom[12] = 120'h00C041D8EC335000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00FA404F8000000000000100113;
    rom[16] = 120'h010300000000000000000000001;
    rom[17] = 120'h0111406E3000000000000120133;
    rom[18] = 120'h012300000000000000000000001;
    rom[19] = 120'h013300000000000000000000001;
    rom[20] = 120'h014A43CA1A63B000000001501C3;
    rom[21] = 120'h015A4360009C400000000160193;
    rom[22] = 120'h0161406E1000000000000170183;
    rom[23] = 120'h017300000000000000000000001;
    rom[24] = 120'h018300000000000000000000000;
    rom[25] = 120'h019041D8EC337000000001A01B3;
    rom[26] = 120'h01A300000000000000000000000;
    rom[27] = 120'h01B300000000000000000000000;
    rom[28] = 120'h01C1407298000000000001D0203;
    rom[29] = 120'h01DA43DF6E4DA000000001E01F3;
    rom[30] = 120'h01E300000000000000000000001;
    rom[31] = 120'h01F300000000000000000000001;
    rom[32] = 120'h020041D8EC33700000000210223;
    rom[33] = 120'h021300000000000000000000000;
    rom[34] = 120'h022300000000000000000000000;
    rom[35] = 120'h0231407388000000000002402D3;
    rom[36] = 120'h024041D8EC337000000002502A3;
    rom[37] = 120'h025140737800000000000260273;
    rom[38] = 120'h026300000000000000000000001;
    rom[39] = 120'h027A405AC000000000000280293;
    rom[40] = 120'h028300000000000000000000000;
    rom[41] = 120'h029300000000000000000000001;
    rom[42] = 120'h02AA414E0ABC0000000002B02C3;
    rom[43] = 120'h02B300000000000000000000000;
    rom[44] = 120'h02C300000000000000000000001;
    rom[45] = 120'h02D300000000000000000000001;
    rom[46] = 120'h02EA4393980AC000000002F04A3;
    rom[47] = 120'h02F041D8EC337000000003003D3;
    rom[48] = 120'h0301407E1800000000000310363;
    rom[49] = 120'h031A4321B60BC00000000320353;
    rom[50] = 120'h032A3FE00000000000000330343;
    rom[51] = 120'h033300000000000000000000000;
    rom[52] = 120'h034300000000000000000000000;
    rom[53] = 120'h035300000000000000000000001;
    rom[54] = 120'h036A432300181000000003703A3;
    rom[55] = 120'h037A40160000000000000380393;
    rom[56] = 120'h038300000000000000000000000;
    rom[57] = 120'h039300000000000000000000000;
    rom[58] = 120'h03A041D8EC335000000003B03C3;
    rom[59] = 120'h03B300000000000000000000001;
    rom[60] = 120'h03C300000000000000000000001;
    rom[61] = 120'h03D1407E18000000000003E0433;
    rom[62] = 120'h03E14077E8000000000003F0403;
    rom[63] = 120'h03F300000000000000000000001;
    rom[64] = 120'h0401407C6800000000000410423;
    rom[65] = 120'h041300000000000000000000000;
    rom[66] = 120'h042300000000000000000000000;
    rom[67] = 120'h043A43230018000000000440473;
    rom[68] = 120'h044A40340000000000000450463;
    rom[69] = 120'h045300000000000000000000000;
    rom[70] = 120'h046300000000000000000000000;
    rom[71] = 120'h047A43250018000000000480493;
    rom[72] = 120'h048300000000000000000000001;
    rom[73] = 120'h049300000000000000000000000;
    rom[74] = 120'h04A041D8EC337000000004B05A3;
    rom[75] = 120'h04BA43D40221F000000004C0533;
    rom[76] = 120'h04CA43B007BB6800000004D0503;
    rom[77] = 120'h04D041D8EC335000000004E04F3;
    rom[78] = 120'h04E300000000000000000000000;
    rom[79] = 120'h04F300000000000000000000000;
    rom[80] = 120'h050140798800000000000510523;
    rom[81] = 120'h051300000000000000000000001;
    rom[82] = 120'h052300000000000000000000000;
    rom[83] = 120'h05314079D800000000000540573;
    rom[84] = 120'h054041D8EC33500000000550563;
    rom[85] = 120'h055300000000000000000000000;
    rom[86] = 120'h056300000000000000000000000;
    rom[87] = 120'h0571407F0800000000000580593;
    rom[88] = 120'h058300000000000000000000001;
    rom[89] = 120'h059300000000000000000000000;
    rom[90] = 120'h05AA43EA5CA1C000000005B0623;
    rom[91] = 120'h05B1407908000000000005C05F3;
    rom[92] = 120'h05C14077D8000000000005D05E3;
    rom[93] = 120'h05D300000000000000000000000;
    rom[94] = 120'h05E300000000000000000000001;
    rom[95] = 120'h05F14079D800000000000600613;
    rom[96] = 120'h060300000000000000000000000;
    rom[97] = 120'h061300000000000000000000000;
    rom[98] = 120'h062300000000000000000000001;
    rom[99] = 120'h0631406BA0000000000006406D3;
    rom[100] = 120'h06414068E000000000000650663;
    rom[101] = 120'h065300000000000000000000000;
    rom[102] = 120'h066A419C00821000000006706C3;
    rom[103] = 120'h067A40C00800000000000680693;
    rom[104] = 120'h068300000000000000000000001;
    rom[105] = 120'h069A418C01042000000006A06B3;
    rom[106] = 120'h06A300000000000000000000000;
    rom[107] = 120'h06B300000000000000000000001;
    rom[108] = 120'h06C300000000000000000000000;
    rom[109] = 120'h06D14075E8000000000006E0773;
    rom[110] = 120'h06E14073C0000000000006F0763;
    rom[111] = 120'h06F1406EA000000000000700713;
    rom[112] = 120'h070300000000000000000000000;
    rom[113] = 120'h07114070C800000000000720753;
    rom[114] = 120'h072041D8EC33B00000000730743;
    rom[115] = 120'h073300000000000000000000000;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h075300000000000000000000000;
    rom[118] = 120'h076300000000000000000000001;
    rom[119] = 120'h077300000000000000000000000;
    rom[120] = 120'h078041D8EC33900000000790BC3;
    rom[121] = 120'h079A3FE000000000000007A08D3;
    rom[122] = 120'h07A041D8EC337000000007B08C3;
    rom[123] = 120'h07B041D8EC335000000007C0853;
    rom[124] = 120'h07C1408880000000000007D07E3;
    rom[125] = 120'h07D300000000000000000000001;
    rom[126] = 120'h07E1409002000000000007F0823;
    rom[127] = 120'h07F1408C5800000000000800813;
    rom[128] = 120'h080300000000000000000000000;
    rom[129] = 120'h081300000000000000000000000;
    rom[130] = 120'h08214092C000000000000830843;
    rom[131] = 120'h083300000000000000000000001;
    rom[132] = 120'h084300000000000000000000000;
    rom[133] = 120'h085140893000000000000860873;
    rom[134] = 120'h086300000000000000000000001;
    rom[135] = 120'h087140918000000000000880893;
    rom[136] = 120'h088300000000000000000000000;
    rom[137] = 120'h08914093B4000000000008A08B3;
    rom[138] = 120'h08A300000000000000000000001;
    rom[139] = 120'h08B300000000000000000000000;
    rom[140] = 120'h08C300000000000000000000000;
    rom[141] = 120'h08DA43A4816EC000000008E0AD3;
    rom[142] = 120'h08E041D8EC337000000008F09E3;
    rom[143] = 120'h08F041D8EC33500000000900973;
    rom[144] = 120'h0901408FDC00000000000910943;
    rom[145] = 120'h091A436FE82AC00000000920933;
    rom[146] = 120'h092300000000000000000000001;
    rom[147] = 120'h093300000000000000000000000;
    rom[148] = 120'h09414093C600000000000950963;
    rom[149] = 120'h095300000000000000000000001;
    rom[150] = 120'h096300000000000000000000001;
    rom[151] = 120'h097A436FE9FD3000000009809B3;
    rom[152] = 120'h098A41701AA87800000009909A3;
    rom[153] = 120'h099300000000000000000000001;
    rom[154] = 120'h09A300000000000000000000001;
    rom[155] = 120'h09B1408E54000000000009C09D3;
    rom[156] = 120'h09C300000000000000000000000;
    rom[157] = 120'h09D300000000000000000000001;
    rom[158] = 120'h09E1408E8C000000000009F0A63;
    rom[159] = 120'h09FA416CFAC8E00000000A00A33;
    rom[160] = 120'h0A01408A3800000000000A10A23;
    rom[161] = 120'h0A1300000000000000000000001;
    rom[162] = 120'h0A2300000000000000000000001;
    rom[163] = 120'h0A31407F5800000000000A40A53;
    rom[164] = 120'h0A4300000000000000000000000;
    rom[165] = 120'h0A5300000000000000000000000;
    rom[166] = 120'h0A6A426C1D38700000000A70AA3;
    rom[167] = 120'h0A71408FCC00000000000A80A93;
    rom[168] = 120'h0A8300000000000000000000001;
    rom[169] = 120'h0A9300000000000000000000001;
    rom[170] = 120'h0AA1408FCC00000000000AB0AC3;
    rom[171] = 120'h0AB300000000000000000000000;
    rom[172] = 120'h0AC300000000000000000000001;
    rom[173] = 120'h0AD14094AA00000000000AE0BB3;
    rom[174] = 120'h0AE1408F4400000000000AF0B63;
    rom[175] = 120'h0AF041D8EC33500000000B00B33;
    rom[176] = 120'h0B0A43AE3BAD500000000B10B23;
    rom[177] = 120'h0B1300000000000000000000000;
    rom[178] = 120'h0B2300000000000000000000001;
    rom[179] = 120'h0B3041D8EC33700000000B40B53;
    rom[180] = 120'h0B4300000000000000000000001;
    rom[181] = 120'h0B5300000000000000000000001;
    rom[182] = 120'h0B6A43E0009EA00000000B70BA3;
    rom[183] = 120'h0B7A43DFFD5F100000000B80B93;
    rom[184] = 120'h0B8300000000000000000000001;
    rom[185] = 120'h0B9300000000000000000000000;
    rom[186] = 120'h0BA300000000000000000000001;
    rom[187] = 120'h0BB300000000000000000000001;
    rom[188] = 120'h0BC041D8EC33B00000000BD0CA3;
    rom[189] = 120'h0BDA421EC808700000000BE0C33;
    rom[190] = 120'h0BEA41E0D730D70000000BF0C03;
    rom[191] = 120'h0BF300000000000000000000000;
    rom[192] = 120'h0C0140890C00000000000C10C23;
    rom[193] = 120'h0C1300000000000000000000000;
    rom[194] = 120'h0C2300000000000000000000001;
    rom[195] = 120'h0C314082E000000000000C40C93;
    rom[196] = 120'h0C4A43A13000080000000C50C63;
    rom[197] = 120'h0C5300000000000000000000000;
    rom[198] = 120'h0C6A43AB1B00000000000C70C83;
    rom[199] = 120'h0C7300000000000000000000001;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C9300000000000000000000000;
    rom[202] = 120'h0CAA43BBF184C00000000CB0D43;
    rom[203] = 120'h0CB1408EE800000000000CC0CD3;
    rom[204] = 120'h0CC300000000000000000000000;
    rom[205] = 120'h0CDA425D680B800000000CE0D33;
    rom[206] = 120'h0CE1408F9000000000000CF0D23;
    rom[207] = 120'h0CFA42140000000000000D00D13;
    rom[208] = 120'h0D0300000000000000000000000;
    rom[209] = 120'h0D1300000000000000000000001;
    rom[210] = 120'h0D2300000000000000000000000;
    rom[211] = 120'h0D3300000000000000000000000;
    rom[212] = 120'h0D4A43BFC403D00000000D50D63;
    rom[213] = 120'h0D5300000000000000000000001;
    rom[214] = 120'h0D6300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 215; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
