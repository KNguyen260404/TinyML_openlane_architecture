module tree_rom_4 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000A43C2154C500000000010CC3;
    rom[1] = 120'h0011408E8C00000000000020873;
    rom[2] = 120'h002041D8EC33900000000030683;
    rom[3] = 120'h003041D8EC33500000000040373;
    rom[4] = 120'h0041406890000000000000501A3;
    rom[5] = 120'h005A436EC661C00000000060113;
    rom[6] = 120'h006A420C2E71B000000000700C3;
    rom[7] = 120'h007A3FE000000000000000800B3;
    rom[8] = 120'h0081405820000000000000900A3;
    rom[9] = 120'h009300000000000000000000001;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00CA42184118D000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E1406810000000000000F0103;
    rom[15] = 120'h00F300000000000000000000001;
    rom[16] = 120'h010300000000000000000000000;
    rom[17] = 120'h011140681000000000000120133;
    rom[18] = 120'h012300000000000000000000001;
    rom[19] = 120'h013A43AC3CED700000000140173;
    rom[20] = 120'h014140683000000000000150163;
    rom[21] = 120'h015300000000000000000000000;
    rom[22] = 120'h016300000000000000000000001;
    rom[23] = 120'h017A43C169D2500000000180193;
    rom[24] = 120'h018300000000000000000000000;
    rom[25] = 120'h019300000000000000000000000;
    rom[26] = 120'h01A1407E58000000000001B02A3;
    rom[27] = 120'h01B14077C8000000000001C0233;
    rom[28] = 120'h01CA435FA1FCB000000001D0203;
    rom[29] = 120'h01DA41DFCE584000000001E01F3;
    rom[30] = 120'h01E300000000000000000000000;
    rom[31] = 120'h01F300000000000000000000001;
    rom[32] = 120'h020A43608BC3800000000210223;
    rom[33] = 120'h021300000000000000000000000;
    rom[34] = 120'h022300000000000000000000000;
    rom[35] = 120'h023A43B1D483500000000240273;
    rom[36] = 120'h024140791800000000000250263;
    rom[37] = 120'h025300000000000000000000000;
    rom[38] = 120'h026300000000000000000000000;
    rom[39] = 120'h027140799800000000000280293;
    rom[40] = 120'h028300000000000000000000001;
    rom[41] = 120'h029300000000000000000000001;
    rom[42] = 120'h02AA3FE000000000000002B0303;
    rom[43] = 120'h02B1408C58000000000002C02F3;
    rom[44] = 120'h02C14088D8000000000002D02E3;
    rom[45] = 120'h02D300000000000000000000000;
    rom[46] = 120'h02E300000000000000000000000;
    rom[47] = 120'h02F300000000000000000000001;
    rom[48] = 120'h030A437003D7200000000310343;
    rom[49] = 120'h031A416A9AF5300000000320333;
    rom[50] = 120'h032300000000000000000000001;
    rom[51] = 120'h033300000000000000000000001;
    rom[52] = 120'h034A43B01A17180000000350363;
    rom[53] = 120'h035300000000000000000000000;
    rom[54] = 120'h036300000000000000000000001;
    rom[55] = 120'h037A43AF83B4300000000380533;
    rom[56] = 120'h038A43A1192AA00000000390483;
    rom[57] = 120'h039041D8EC337000000003A0413;
    rom[58] = 120'h03AA4374A80AB000000003B03E3;
    rom[59] = 120'h03B1406810000000000003C03D3;
    rom[60] = 120'h03C300000000000000000000001;
    rom[61] = 120'h03D300000000000000000000000;
    rom[62] = 120'h03EA439925C4A000000003F0403;
    rom[63] = 120'h03F300000000000000000000000;
    rom[64] = 120'h040300000000000000000000000;
    rom[65] = 120'h0411406E1000000000000420453;
    rom[66] = 120'h042A42F4B75A700000000430443;
    rom[67] = 120'h043300000000000000000000001;
    rom[68] = 120'h044300000000000000000000000;
    rom[69] = 120'h045A43229F79800000000460473;
    rom[70] = 120'h046300000000000000000000000;
    rom[71] = 120'h047300000000000000000000000;
    rom[72] = 120'h0481407E98000000000004904E3;
    rom[73] = 120'h0491407E48000000000004A04B3;
    rom[74] = 120'h04A300000000000000000000001;
    rom[75] = 120'h04BA43AD516F2000000004C04D3;
    rom[76] = 120'h04C300000000000000000000001;
    rom[77] = 120'h04D300000000000000000000000;
    rom[78] = 120'h04EA43AE1D4E3000000004F0503;
    rom[79] = 120'h04F300000000000000000000001;
    rom[80] = 120'h050041D8EC33700000000510523;
    rom[81] = 120'h051300000000000000000000000;
    rom[82] = 120'h052300000000000000000000001;
    rom[83] = 120'h053A43B0E043F000000005405B3;
    rom[84] = 120'h0541407F18000000000005505A3;
    rom[85] = 120'h055140669000000000000560573;
    rom[86] = 120'h056300000000000000000000001;
    rom[87] = 120'h057A43B068D7C00000000580593;
    rom[88] = 120'h058300000000000000000000000;
    rom[89] = 120'h059300000000000000000000000;
    rom[90] = 120'h05A300000000000000000000001;
    rom[91] = 120'h05B14068B0000000000005C0613;
    rom[92] = 120'h05C1406810000000000005D05E3;
    rom[93] = 120'h05D300000000000000000000001;
    rom[94] = 120'h05E1406890000000000005F0603;
    rom[95] = 120'h05F300000000000000000000000;
    rom[96] = 120'h060300000000000000000000000;
    rom[97] = 120'h061041D8EC33700000000620653;
    rom[98] = 120'h062A43C1FD0DE00000000630643;
    rom[99] = 120'h063300000000000000000000001;
    rom[100] = 120'h064300000000000000000000001;
    rom[101] = 120'h0651407F6800000000000660673;
    rom[102] = 120'h066300000000000000000000001;
    rom[103] = 120'h067300000000000000000000001;
    rom[104] = 120'h068041D8EC33B00000000690863;
    rom[105] = 120'h069A419C00821000000006A0753;
    rom[106] = 120'h06AA403300000000000006B06C3;
    rom[107] = 120'h06B300000000000000000000000;
    rom[108] = 120'h06CA405680000000000006D06E3;
    rom[109] = 120'h06D300000000000000000000001;
    rom[110] = 120'h06E1406BA0000000000006F0723;
    rom[111] = 120'h06FA418C0104200000000700713;
    rom[112] = 120'h070300000000000000000000000;
    rom[113] = 120'h071300000000000000000000001;
    rom[114] = 120'h072A41300104800000000730743;
    rom[115] = 120'h073300000000000000000000000;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h075A42D000002000000007607F3;
    rom[118] = 120'h07614070C8000000000007707A3;
    rom[119] = 120'h0771406EA000000000000780793;
    rom[120] = 120'h078300000000000000000000000;
    rom[121] = 120'h079300000000000000000000001;
    rom[122] = 120'h07A1408A48000000000007B07C3;
    rom[123] = 120'h07B300000000000000000000000;
    rom[124] = 120'h07CA4201C1B515C0000007D07E3;
    rom[125] = 120'h07D300000000000000000000000;
    rom[126] = 120'h07E300000000000000000000001;
    rom[127] = 120'h07F1407EF000000000000800813;
    rom[128] = 120'h080300000000000000000000000;
    rom[129] = 120'h08114086D800000000000820853;
    rom[130] = 120'h082A43A13000080000000830843;
    rom[131] = 120'h083300000000000000000000000;
    rom[132] = 120'h084300000000000000000000000;
    rom[133] = 120'h085300000000000000000000000;
    rom[134] = 120'h086300000000000000000000000;
    rom[135] = 120'h087A3FE000000000000008809B3;
    rom[136] = 120'h08814099F0000000000008909A3;
    rom[137] = 120'h089041D8EC337000000008A0993;
    rom[138] = 120'h08A041D8EC335000000008B0923;
    rom[139] = 120'h08B140950C000000000008C0913;
    rom[140] = 120'h08C1409002000000000008D08E3;
    rom[141] = 120'h08D300000000000000000000000;
    rom[142] = 120'h08E14092C0000000000008F0903;
    rom[143] = 120'h08F300000000000000000000001;
    rom[144] = 120'h090300000000000000000000000;
    rom[145] = 120'h091300000000000000000000001;
    rom[146] = 120'h092140943600000000000930983;
    rom[147] = 120'h09314091AA00000000000940953;
    rom[148] = 120'h094300000000000000000000000;
    rom[149] = 120'h09514093B4000000000001200973;
    rom[150] = 120'h0120300000000000000000000001;
    rom[151] = 120'h097300000000000000000000000;
    rom[152] = 120'h098300000000000000000000001;
    rom[153] = 120'h099300000000000000000000000;
    rom[154] = 120'h09A300000000000000000000000;
    rom[155] = 120'h09B041D8EC33B000000009C0BF3;
    rom[156] = 120'h09CA426C2589E000000009D0AE3;
    rom[157] = 120'h09D041D8EC339000000009E0AB3;
    rom[158] = 120'h09EA408404000000000009F0A43;
    rom[159] = 120'h09F1408FE000000000000A00A33;
    rom[160] = 120'h0A0041D8EC33700000000A10A23;
    rom[161] = 120'h0A1300000000000000000000000;
    rom[162] = 120'h0A2300000000000000000000000;
    rom[163] = 120'h0A3300000000000000000000001;
    rom[164] = 120'h0A4041D8EC33500000000A50A83;
    rom[165] = 120'h0A5A41D67BC6400000000A60A73;
    rom[166] = 120'h0A6300000000000000000000001;
    rom[167] = 120'h0A7300000000000000000000001;
    rom[168] = 120'h0A8041D8EC33700000000A90AA3;
    rom[169] = 120'h0A9300000000000000000000001;
    rom[170] = 120'h0AA300000000000000000000001;
    rom[171] = 120'h0AB1408F9000000000000AC0AD3;
    rom[172] = 120'h0AC300000000000000000000001;
    rom[173] = 120'h0AD300000000000000000000000;
    rom[174] = 120'h0AE041D8EC33900000000AF0BE3;
    rom[175] = 120'h0AF041D8EC33500000000B00B73;
    rom[176] = 120'h0B01408FCC00000000000B10B43;
    rom[177] = 120'h0B1A42F04B84A00000000B20B33;
    rom[178] = 120'h0B2300000000000000000000001;
    rom[179] = 120'h0B3300000000000000000000000;
    rom[180] = 120'h0B4A426C2A2C200000000B50B63;
    rom[181] = 120'h0B5300000000000000000000000;
    rom[182] = 120'h0B6300000000000000000000001;
    rom[183] = 120'h0B7041D8EC33700000000B80BB3;
    rom[184] = 120'h0B8A43C21136F00000000B90BA3;
    rom[185] = 120'h0B9300000000000000000000001;
    rom[186] = 120'h0BA300000000000000000000000;
    rom[187] = 120'h0BBA43B33B1C200000000BC0BD3;
    rom[188] = 120'h0BC300000000000000000000000;
    rom[189] = 120'h0BD300000000000000000000001;
    rom[190] = 120'h0BE300000000000000000000000;
    rom[191] = 120'h0BF041D8EC33D00000000C00C53;
    rom[192] = 120'h0C0A43BBEF84800000000C10C23;
    rom[193] = 120'h0C1300000000000000000000000;
    rom[194] = 120'h0C2A43C02A4F380000000C30C43;
    rom[195] = 120'h0C3300000000000000000000001;
    rom[196] = 120'h0C4300000000000000000000000;
    rom[197] = 120'h0C51408F6800000000000C60CB3;
    rom[198] = 120'h0C6041D8EC33F00000000C70CA3;
    rom[199] = 120'h0C7A42A22800000000000C80C93;
    rom[200] = 120'h0C8300000000000000000000001;
    rom[201] = 120'h0C9300000000000000000000000;
    rom[202] = 120'h0CA300000000000000000000000;
    rom[203] = 120'h0CB300000000000000000000000;
    rom[204] = 120'h0CC140681000000000000CD0CE3;
    rom[205] = 120'h0CD300000000000000000000001;
    rom[206] = 120'h0CEA43D3FFE4D00000000CF0F63;
    rom[207] = 120'h0CF1407F5800000000000D00E93;
    rom[208] = 120'h0D01407E9800000000000D10E03;
    rom[209] = 120'h0D1041D8EC33900000000D20DF3;
    rom[210] = 120'h0D2041D8EC33700000000D30DA3;
    rom[211] = 120'h0D31407E4800000000000D40D73;
    rom[212] = 120'h0D4A43C7FFB4800000000D50D63;
    rom[213] = 120'h0D5300000000000000000000001;
    rom[214] = 120'h0D6300000000000000000000000;
    rom[215] = 120'h0D7041D8EC33500000000D80D93;
    rom[216] = 120'h0D8300000000000000000000000;
    rom[217] = 120'h0D9300000000000000000000000;
    rom[218] = 120'h0DAA43C7BE9F500000000DB0DC3;
    rom[219] = 120'h0DB300000000000000000000001;
    rom[220] = 120'h0DC140797000000000000DD0DE3;
    rom[221] = 120'h0DD300000000000000000000000;
    rom[222] = 120'h0DE300000000000000000000000;
    rom[223] = 120'h0DF300000000000000000000000;
    rom[224] = 120'h0E01407F4800000000000E10E23;
    rom[225] = 120'h0E1300000000000000000000001;
    rom[226] = 120'h0E2A43D14340000000000E30E83;
    rom[227] = 120'h0E3041D8EC33500000000E40E53;
    rom[228] = 120'h0E4300000000000000000000001;
    rom[229] = 120'h0E5041D8EC33700000000E60E73;
    rom[230] = 120'h0E6300000000000000000000000;
    rom[231] = 120'h0E7300000000000000000000000;
    rom[232] = 120'h0E8300000000000000000000001;
    rom[233] = 120'h0E9140932200000000000EA0EB3;
    rom[234] = 120'h0EA300000000000000000000001;
    rom[235] = 120'h0EBA43D007FE700000000EC0ED3;
    rom[236] = 120'h0EC300000000000000000000001;
    rom[237] = 120'h0ED140945200000000000EE0F53;
    rom[238] = 120'h0EE041D8EC33700000000EF0F23;
    rom[239] = 120'h0EFA43D1D2B3E00000000F00F13;
    rom[240] = 120'h0F0300000000000000000000000;
    rom[241] = 120'h0F1300000000000000000000001;
    rom[242] = 120'h0F2041D8EC33900000000F30F43;
    rom[243] = 120'h0F3300000000000000000000000;
    rom[244] = 120'h0F4300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 

