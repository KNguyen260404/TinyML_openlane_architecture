module tree_rom_5 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000140681000000000000010023;
    rom[1] = 120'h001300000000000000000000001;
    rom[2] = 120'h0021407F38000000000000306C3;
    rom[3] = 120'h00314077C8000000000000403D3;
    rom[4] = 120'h004140734800000000000050303;
    rom[5] = 120'h0051406E1000000000000060213;
    rom[6] = 120'h006A43600097B00000000070143;
    rom[7] = 120'h0071406890000000000000800F3;
    rom[8] = 120'h008041D8EC335000000000900C3;
    rom[9] = 120'h009A4203FB67E000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000000;
    rom[12] = 120'h00C1406830000000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00F041D8EC33B00000000100133;
    rom[16] = 120'h010041D8EC33500000000110123;
    rom[17] = 120'h011300000000000000000000001;
    rom[18] = 120'h012300000000000000000000001;
    rom[19] = 120'h013300000000000000000000000;
    rom[20] = 120'h014041D8EC337000000001501C3;
    rom[21] = 120'h015041D8EC33500000000160193;
    rom[22] = 120'h016140693000000000000170183;
    rom[23] = 120'h017300000000000000000000000;
    rom[24] = 120'h018300000000000000000000001;
    rom[25] = 120'h019A43CA2830F000000001A01B3;
    rom[26] = 120'h01A300000000000000000000000;
    rom[27] = 120'h01B300000000000000000000001;
    rom[28] = 120'h01C041D8EC339000000001D0203;
    rom[29] = 120'h01DA43CA4043F000000001E01F3;
    rom[30] = 120'h01E300000000000000000000000;
    rom[31] = 120'h01F300000000000000000000001;
    rom[32] = 120'h020300000000000000000000000;
    rom[33] = 120'h021A43DF81ECE000000002202F3;
    rom[34] = 120'h022A40AFDC00000000000230283;
    rom[35] = 120'h023A40502000000000000240273;
    rom[36] = 120'h0241406E3000000000000250263;
    rom[37] = 120'h025300000000000000000000000;
    rom[38] = 120'h026300000000000000000000001;
    rom[39] = 120'h027300000000000000000000001;
    rom[40] = 120'h0281406F30000000000002902C3;
    rom[41] = 120'h0291406E30000000000002A02B3;
    rom[42] = 120'h02A300000000000000000000000;
    rom[43] = 120'h02B300000000000000000000000;
    rom[44] = 120'h02C041D8EC337000000002D02E3;
    rom[45] = 120'h02D300000000000000000000001;
    rom[46] = 120'h02E300000000000000000000000;
    rom[47] = 120'h02F300000000000000000000001;
    rom[48] = 120'h030041D8EC33B000000003103C3;
    rom[49] = 120'h031041D8EC33900000000320393;
    rom[50] = 120'h032140738800000000000330383;
    rom[51] = 120'h033140737800000000000340353;
    rom[52] = 120'h034300000000000000000000001;
    rom[53] = 120'h035A403E8000000000000360373;
    rom[54] = 120'h036300000000000000000000000;
    rom[55] = 120'h037300000000000000000000001;
    rom[56] = 120'h038300000000000000000000001;
    rom[57] = 120'h039A412002140000000003A03B3;
    rom[58] = 120'h03A300000000000000000000000;
    rom[59] = 120'h03B300000000000000000000001;
    rom[60] = 120'h03C300000000000000000000000;
    rom[61] = 120'h03D041D8EC339000000003E06B3;
    rom[62] = 120'h03E1407E58000000000003F0543;
    rom[63] = 120'h03F1407E08000000000004004D3;
    rom[64] = 120'h040041D8EC33700000000410483;
    rom[65] = 120'h041041D8EC33500000000420453;
    rom[66] = 120'h0421407CD800000000000430443;
    rom[67] = 120'h043300000000000000000000000;
    rom[68] = 120'h044300000000000000000000001;
    rom[69] = 120'h0451407CD800000000000460473;
    rom[70] = 120'h046300000000000000000000000;
    rom[71] = 120'h047300000000000000000000001;
    rom[72] = 120'h048A43EA18721000000004904C3;
    rom[73] = 120'h049A43B0B07F1000000004A04B3;
    rom[74] = 120'h04A300000000000000000000000;
    rom[75] = 120'h04B300000000000000000000000;
    rom[76] = 120'h04C300000000000000000000001;
    rom[77] = 120'h04DA43D1DEB76000000004E0533;
    rom[78] = 120'h04EA4120F7AF0000000004F0503;
    rom[79] = 120'h04F300000000000000000000001;
    rom[80] = 120'h0501407E4800000000000510523;
    rom[81] = 120'h051300000000000000000000000;
    rom[82] = 120'h052300000000000000000000000;
    rom[83] = 120'h053300000000000000000000001;
    rom[84] = 120'h054A43240018100000000550623;
    rom[85] = 120'h055A432300181000000005605B3;
    rom[86] = 120'h0561407E8800000000000570583;
    rom[87] = 120'h057300000000000000000000001;
    rom[88] = 120'h0581407F28000000000005905A3;
    rom[89] = 120'h059300000000000000000000000;
    rom[90] = 120'h05A300000000000000000000000;
    rom[91] = 120'h05B041D8EC335000000005C05F3;
    rom[92] = 120'h05C1407EA0000000000005D05E3;
    rom[93] = 120'h05D300000000000000000000001;
    rom[94] = 120'h05E300000000000000000000001;
    rom[95] = 120'h05F041D8EC33700000000600613;
    rom[96] = 120'h060300000000000000000000001;
    rom[97] = 120'h061300000000000000000000001;
    rom[98] = 120'h0621407E8800000000000630643;
    rom[99] = 120'h063300000000000000000000001;
    rom[100] = 120'h064041D8EC33500000000650683;
    rom[101] = 120'h0651407E9800000000000660673;
    rom[102] = 120'h066300000000000000000000000;
    rom[103] = 120'h067300000000000000000000000;
    rom[104] = 120'h068041D8EC337000000006906A3;
    rom[105] = 120'h069300000000000000000000000;
    rom[106] = 120'h06A300000000000000000000000;
    rom[107] = 120'h06B300000000000000000000000;
    rom[108] = 120'h06C041D8EC339000000006D0C03;
    rom[109] = 120'h06D1408FDC000000000006E0993;
    rom[110] = 120'h06E041D8EC337000000006F0803;
    rom[111] = 120'h06FA3FE00000000000000700733;
    rom[112] = 120'h07014088D400000000000710723;
    rom[113] = 120'h071300000000000000000000001;
    rom[114] = 120'h072300000000000000000000000;
    rom[115] = 120'h0731408F64000000000007407B3;
    rom[116] = 120'h074041D8EC33500000000750783;
    rom[117] = 120'h0751407F5800000000000760773;
    rom[118] = 120'h076300000000000000000000000;
    rom[119] = 120'h077300000000000000000000001;
    rom[120] = 120'h0781408614000000000007907A3;
    rom[121] = 120'h079300000000000000000000001;
    rom[122] = 120'h07A300000000000000000000001;
    rom[123] = 120'h07BA43E000904000000007C07F3;
    rom[124] = 120'h07C041D8EC335000000007D07E3;
    rom[125] = 120'h07D300000000000000000000000;
    rom[126] = 120'h07E300000000000000000000000;
    rom[127] = 120'h07F300000000000000000000001;
    rom[128] = 120'h0801408614000000000008108C3;
    rom[129] = 120'h081A4391C380800000000820873;
    rom[130] = 120'h0821407F5800000000000830863;
    rom[131] = 120'h0831407F4800000000000840853;
    rom[132] = 120'h084300000000000000000000001;
    rom[133] = 120'h085300000000000000000000000;
    rom[134] = 120'h086300000000000000000000001;
    rom[135] = 120'h0871407F58000000000008808B3;
    rom[136] = 120'h088A43C16E135000000008908A3;
    rom[137] = 120'h089300000000000000000000001;
    rom[138] = 120'h08A300000000000000000000000;
    rom[139] = 120'h08B300000000000000000000001;
    rom[140] = 120'h08CA41AAE460C000000008D0923;
    rom[141] = 120'h08DA3FF000000000000008E08F3;
    rom[142] = 120'h08E300000000000000000000000;
    rom[143] = 120'h08FA416ECAA6900000000900913;
    rom[144] = 120'h090300000000000000000000001;
    rom[145] = 120'h091300000000000000000000000;
    rom[146] = 120'h0921408E8C000000000009301203;
    rom[147] = 120'h0931408E0400000000000940953;
    rom[148] = 120'h094300000000000000000000000;
    rom[149] = 120'h095300000000000000000000000;
    rom[150] = 120'h0120A43DF7498A00000000970983;
    rom[151] = 120'h097300000000000000000000001;
    rom[152] = 120'h098300000000000000000000000;
    rom[153] = 120'h099041D8EC337000000009A0B33;
    rom[154] = 120'h09A14094AA000000000009B0A83;
    rom[155] = 120'h09BA3FE000000000000009C0A13;
    rom[156] = 120'h09C14093B4000000000009D09E3;
    rom[157] = 120'h09D300000000000000000000001;
    rom[158] = 120'h09E1409436000000000009F0A03;
    rom[159] = 120'h09F300000000000000000000000;
    rom[160] = 120'h0A0300000000000000000000001;
    rom[161] = 120'h0A1041D8EC33500000000A20A53;
    rom[162] = 120'h0A2A43D1CCAD000000000A30A43;
    rom[163] = 120'h0A3300000000000000000000001;
    rom[164] = 120'h0A4300000000000000000000001;
    rom[165] = 120'h0A5A43D1DAB3300000000A60A73;
    rom[166] = 120'h0A6300000000000000000000001;
    rom[167] = 120'h0A7300000000000000000000001;
    rom[168] = 120'h0A8A3FE00000000000000A90AE3;
    rom[169] = 120'h0A9041D8EC33500000000AA0AD3;
    rom[170] = 120'h0AA1409D5E00000000000AB0AC3;
    rom[171] = 120'h0AB300000000000000000000001;
    rom[172] = 120'h0AC300000000000000000000000;
    rom[173] = 120'h0AD300000000000000000000000;
    rom[174] = 120'h0AE1409DC200000000000AF0B03;
    rom[175] = 120'h0AF300000000000000000000001;
    rom[176] = 120'h0B01409DCE00000000000B10B23;
    rom[177] = 120'h0B1300000000000000000000001;
    rom[178] = 120'h0B2300000000000000000000001;
    rom[179] = 120'h0B3A3FF00000000000000B40B53;
    rom[180] = 120'h0B4300000000000000000000000;
    rom[181] = 120'h0B514094AC00000000000B60BB3;
    rom[182] = 120'h0B6A426C1D38700000000B70B83;
    rom[183] = 120'h0B7300000000000000000000001;
    rom[184] = 120'h0B8A43D1CC72B00000000B90BA3;
    rom[185] = 120'h0B9300000000000000000000000;
    rom[186] = 120'h0BA300000000000000000000001;
    rom[187] = 120'h0BB1409DC200000000000BC0BD3;
    rom[188] = 120'h0BC300000000000000000000001;
    rom[189] = 120'h0BDA42D40713900000000BE0BF3;
    rom[190] = 120'h0BE300000000000000000000001;
    rom[191] = 120'h0BF300000000000000000000001;
    rom[192] = 120'h0C0041D8EC33B00000000C10CE3;
    rom[193] = 120'h0C1A421EC808700000000C20C73;
    rom[194] = 120'h0C2A41E0D730D70000000C30C43;
    rom[195] = 120'h0C3300000000000000000000000;
    rom[196] = 120'h0C4140890C00000000000C50C63;
    rom[197] = 120'h0C5300000000000000000000000;
    rom[198] = 120'h0C6300000000000000000000001;
    rom[199] = 120'h0C7A43A9D717D00000000C80C93;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C9140877800000000000CA0CD3;
    rom[202] = 120'h0CAA43AB1B00000000000CB0CC3;
    rom[203] = 120'h0CB300000000000000000000001;
    rom[204] = 120'h0CC300000000000000000000000;
    rom[205] = 120'h0CD300000000000000000000000;
    rom[206] = 120'h0CE041D8EC33D00000000CF0D63;
    rom[207] = 120'h0CFA43BBF184C00000000D00D13;
    rom[208] = 120'h0D0300000000000000000000000;
    rom[209] = 120'h0D11408F5800000000000D20D53;
    rom[210] = 120'h0D2140877800000000000D30D43;
    rom[211] = 120'h0D3300000000000000000000000;
    rom[212] = 120'h0D4300000000000000000000001;
    rom[213] = 120'h0D5300000000000000000000000;
    rom[214] = 120'h0D61408EE800000000000D70D83;
    rom[215] = 120'h0D7300000000000000000000000;
    rom[216] = 120'h0D81408F5800000000000D90DE3;
    rom[217] = 120'h0D9A42A05800000000000DA0DD3;
    rom[218] = 120'h0DAA42140000000000000DB0DC3;
    rom[219] = 120'h0DB300000000000000000000000;
    rom[220] = 120'h0DC300000000000000000000001;
    rom[221] = 120'h0DD300000000000000000000000;
    rom[222] = 120'h0DE300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 223; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 

