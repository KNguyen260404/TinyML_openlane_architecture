module tree_rom_11 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000A43C2154C500000000010B23;
    rom[1] = 120'h0011408E8C00000000000020793;
    rom[2] = 120'h002041D8EC339000000000305A3;
    rom[3] = 120'h003140689000000000000040293;
    rom[4] = 120'h004A436D5F10D00000000050143;
    rom[5] = 120'h005A420F94B9F000000000600D3;
    rom[6] = 120'h006A3FE000000000000000700C3;
    rom[7] = 120'h00714066B000000000000080093;
    rom[8] = 120'h008300000000000000000000001;
    rom[9] = 120'h009041D8EC335000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000000;
    rom[12] = 120'h00C300000000000000000000001;
    rom[13] = 120'h00D1406810000000000000E00F3;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00F140683000000000000100133;
    rom[16] = 120'h010041D8EC33500000000110123;
    rom[17] = 120'h011300000000000000000000000;
    rom[18] = 120'h012300000000000000000000000;
    rom[19] = 120'h013300000000000000000000001;
    rom[20] = 120'h014A43BFF8BCB00000000150203;
    rom[21] = 120'h015A43B40343E000000001601B3;
    rom[22] = 120'h016140681000000000000170183;
    rom[23] = 120'h017300000000000000000000001;
    rom[24] = 120'h0181406830000000000001901A3;
    rom[25] = 120'h019300000000000000000000000;
    rom[26] = 120'h01A300000000000000000000001;
    rom[27] = 120'h01B041D8EC335000000001C01F3;
    rom[28] = 120'h01CA43B818EB1000000001D01E3;
    rom[29] = 120'h01D300000000000000000000001;
    rom[30] = 120'h01E300000000000000000000001;
    rom[31] = 120'h01F300000000000000000000001;
    rom[32] = 120'h020A43C1FFFD500000000210283;
    rom[33] = 120'h021A43C0210E700000000220253;
    rom[34] = 120'h022140667000000000000230243;
    rom[35] = 120'h023300000000000000000000001;
    rom[36] = 120'h024300000000000000000000000;
    rom[37] = 120'h02514067E000000000000260273;
    rom[38] = 120'h026300000000000000000000001;
    rom[39] = 120'h027300000000000000000000000;
    rom[40] = 120'h028300000000000000000000001;
    rom[41] = 120'h029A400400000000000002A03B3;
    rom[42] = 120'h02A14076F8000000000002B0303;
    rom[43] = 120'h02BA3FF800000000000002C02F3;
    rom[44] = 120'h02C1406920000000000002D02E3;
    rom[45] = 120'h02D300000000000000000000000;
    rom[46] = 120'h02E300000000000000000000001;
    rom[47] = 120'h02F300000000000000000000000;
    rom[48] = 120'h030041D8EC33500000000310363;
    rom[49] = 120'h0311408C5800000000000320353;
    rom[50] = 120'h032A3FE00000000000000330343;
    rom[51] = 120'h033300000000000000000000000;
    rom[52] = 120'h034300000000000000000000001;
    rom[53] = 120'h035300000000000000000000001;
    rom[54] = 120'h036A3FE000000000000003703A3;
    rom[55] = 120'h037041D8EC33700000000380393;
    rom[56] = 120'h038300000000000000000000000;
    rom[57] = 120'h039300000000000000000000000;
    rom[58] = 120'h03A300000000000000000000001;
    rom[59] = 120'h03BA40F001780000000003C04B3;
    rom[60] = 120'h03CA406FD0000000000003D0443;
    rom[61] = 120'h03DA404F40000000000003E0413;
    rom[62] = 120'h03E041D8EC335000000003F0403;
    rom[63] = 120'h03F300000000000000000000001;
    rom[64] = 120'h040300000000000000000000001;
    rom[65] = 120'h041A40502000000000000420433;
    rom[66] = 120'h042300000000000000000000000;
    rom[67] = 120'h043300000000000000000000001;
    rom[68] = 120'h044041D8EC33700000000450483;
    rom[69] = 120'h045A40B01580000000000460473;
    rom[70] = 120'h046300000000000000000000000;
    rom[71] = 120'h047300000000000000000000001;
    rom[72] = 120'h04814079E8000000000004904A3;
    rom[73] = 120'h049300000000000000000000000;
    rom[74] = 120'h04A300000000000000000000001;
    rom[75] = 120'h04B1407E58000000000004C0533;
    rom[76] = 120'h04C041D8EC337000000004D0503;
    rom[77] = 120'h04D14077C8000000000004E04F3;
    rom[78] = 120'h04E300000000000000000000000;
    rom[79] = 120'h04F300000000000000000000000;
    rom[80] = 120'h05014077C800000000000510523;
    rom[81] = 120'h051300000000000000000000000;
    rom[82] = 120'h052300000000000000000000000;
    rom[83] = 120'h053A42A26B7A100000000540573;
    rom[84] = 120'h054A416FFF67C00000000550563;
    rom[85] = 120'h055300000000000000000000001;
    rom[86] = 120'h056300000000000000000000000;
    rom[87] = 120'h057A43240018100000000580593;
    rom[88] = 120'h058300000000000000000000001;
    rom[89] = 120'h059300000000000000000000001;
    rom[90] = 120'h05A1406BA0000000000005B0663;
    rom[91] = 120'h05B14068E0000000000005C05D3;
    rom[92] = 120'h05C300000000000000000000000;
    rom[93] = 120'h05D041D8EC33B000000005E0653;
    rom[94] = 120'h05EA419C00821000000005F0643;
    rom[95] = 120'h05FA40C00800000000000600613;
    rom[96] = 120'h060300000000000000000000001;
    rom[97] = 120'h061A418C0104200000000620633;
    rom[98] = 120'h062300000000000000000000000;
    rom[99] = 120'h063300000000000000000000001;
    rom[100] = 120'h064300000000000000000000000;
    rom[101] = 120'h065300000000000000000000000;
    rom[102] = 120'h06614075E800000000000670703;
    rom[103] = 120'h06714073C0000000000006806F3;
    rom[104] = 120'h0681406EA0000000000006906A3;
    rom[105] = 120'h069300000000000000000000000;
    rom[106] = 120'h06A14070C8000000000006B06E3;
    rom[107] = 120'h06B041D8EC33B000000006C06D3;
    rom[108] = 120'h06C300000000000000000000000;
    rom[109] = 120'h06D300000000000000000000000;
    rom[110] = 120'h06E300000000000000000000000;
    rom[111] = 120'h06F300000000000000000000001;
    rom[112] = 120'h070A420D9010E00000000710723;
    rom[113] = 120'h071300000000000000000000000;
    rom[114] = 120'h072A421EC608700000000730743;
    rom[115] = 120'h073300000000000000000000001;
    rom[116] = 120'h074A43A56208500000000750763;
    rom[117] = 120'h075300000000000000000000000;
    rom[118] = 120'h076041D8EC33B00000000770783;
    rom[119] = 120'h077300000000000000000000000;
    rom[120] = 120'h078300000000000000000000000;
    rom[121] = 120'h079041D8EC33B000000007A0A73;
    rom[122] = 120'h07A041D8EC339000000007B0A23;
    rom[123] = 120'h07BA3FE000000000000007C0853;
    rom[124] = 120'h07C041D8EC337000000007D0843;
    rom[125] = 120'h07D14090B6000000000007E07F3;
    rom[126] = 120'h07E300000000000000000000000;
    rom[127] = 120'h07F14093B400000000000800813;
    rom[128] = 120'h080300000000000000000000001;
    rom[129] = 120'h0811409D5E00000000000820833;
    rom[130] = 120'h082300000000000000000000000;
    rom[131] = 120'h083300000000000000000000000;
    rom[132] = 120'h084300000000000000000000000;
    rom[133] = 120'h085A426C2450F00000000860933;
    rom[134] = 120'h086A40838C000000000008708C3;
    rom[135] = 120'h0871408FE4000000000008808B3;
    rom[136] = 120'h088041D8EC337000000008908A3;
    rom[137] = 120'h089300000000000000000000000;
    rom[138] = 120'h08A300000000000000000000000;
    rom[139] = 120'h08B300000000000000000000001;
    rom[140] = 120'h08C041D8EC335000000008D0903;
    rom[141] = 120'h08D1408FCC000000000008E08F3;
    rom[142] = 120'h08E300000000000000000000001;
    rom[143] = 120'h08F300000000000000000000001;
    rom[144] = 120'h0901408FCC00000000000910923;
    rom[145] = 120'h091300000000000000000000001;
    rom[146] = 120'h092300000000000000000000001;
    rom[147] = 120'h09314093C6000000000009409B3;
    rom[148] = 120'h094041D8EC33700000000950983;
    rom[149] = 120'h095A4367C4D3F00000000960973;
    rom[150] = 120'h096300000000000000000000001;
    rom[151] = 120'h097300000000000000000000001;
    rom[152] = 120'h0981408F80000000000009909A3;
    rom[153] = 120'h099300000000000000000000001;
    rom[154] = 120'h09A300000000000000000000000;
    rom[155] = 120'h09B041D8EC337000000009C09F3;
    rom[156] = 120'h09CA43C20FEBF000000009D09E3;
    rom[157] = 120'h09D300000000000000000000001;
    rom[158] = 120'h09E300000000000000000000000;
    rom[159] = 120'h09FA42D01124400000000A00A13;
    rom[160] = 120'h0A0300000000000000000000001;
    rom[161] = 120'h0A1300000000000000000000001;
    rom[162] = 120'h0A21408F6800000000000A30A63;
    rom[163] = 120'h0A3A42651000400000000A40A53;
    rom[164] = 120'h0A4300000000000000000000001;
    rom[165] = 120'h0A5300000000000000000000000;
    rom[166] = 120'h0A6300000000000000000000000;
    rom[167] = 120'h0A7041D8EC33D00000000A80AD3;
    rom[168] = 120'h0A8A43BBF184C00000000A90AA3;
    rom[169] = 120'h0A9300000000000000000000000;
    rom[170] = 120'h0AA140922600000000000AB0AC3;
    rom[171] = 120'h0AB300000000000000000000001;
    rom[172] = 120'h0AC300000000000000000000000;
    rom[173] = 120'h0ADA425D680B800000000AE0B13;
    rom[174] = 120'h0AEA42140000040000000AF0B03;
    rom[175] = 120'h0AF300000000000000000000000;
    rom[176] = 120'h0B0300000000000000000000001;
    rom[177] = 120'h0B1300000000000000000000000;
    rom[178] = 120'h0B2A43C7FFB4800000000B30B43;
    rom[179] = 120'h0B3300000000000000000000001;
    rom[180] = 120'h0B41407F5800000000000B50F63;
    rom[181] = 120'h0B5140798800000000000B60D13;
    rom[182] = 120'h0B6A43D1C0F4C00000000B70C63;
    rom[183] = 120'h0B7041D8EC33900000000B80C53;
    rom[184] = 120'h0B8A43CA0754300000000B90BE3;
    rom[185] = 120'h0B9A43C80412200000000BA0BB3;
    rom[186] = 120'h0BA300000000000000000000000;
    rom[187] = 120'h0BBA43C8042F100000000BC0BD3;
    rom[188] = 120'h0BC300000000000000000000001;
    rom[189] = 120'h0BD300000000000000000000000;
    rom[190] = 120'h0BE140729800000000000BF0C23;
    rom[191] = 120'h0BF140683000000000000C00C13;
    rom[192] = 120'h0C0300000000000000000000001;
    rom[193] = 120'h0C1300000000000000000000001;
    rom[194] = 120'h0C2A43D1B8BB300000000C30C43;
    rom[195] = 120'h0C3300000000000000000000001;
    rom[196] = 120'h0C4300000000000000000000000;
    rom[197] = 120'h0C5300000000000000000000000;
    rom[198] = 120'h0C6A43DED856400000000C70C83;
    rom[199] = 120'h0C7300000000000000000000001;
    rom[200] = 120'h0C81406F1000000000000C90CA3;
    rom[201] = 120'h0C9300000000000000000000001;
    rom[202] = 120'h0CA041D8EC33500000000CB0CE3;
    rom[203] = 120'h0CB1406F3000000000000CC0CD3;
    rom[204] = 120'h0CC300000000000000000000000;
    rom[205] = 120'h0CD300000000000000000000001;
    rom[206] = 120'h0CEA43DF4C99300000000CF0D03;
    rom[207] = 120'h0CF300000000000000000000000;
    rom[208] = 120'h0D0300000000000000000000001;
    rom[209] = 120'h0D1A43EA3A6F100000000D20EB3;
    rom[210] = 120'h0D2041D8EC33700000000D30E03;
    rom[211] = 120'h0D31407F1800000000000D40DB3;
    rom[212] = 120'h0D414079D800000000000D50D83;
    rom[213] = 120'h0D5041D8EC33500000000D60D73;
    rom[214] = 120'h0D6300000000000000000000000;
    rom[215] = 120'h0D7300000000000000000000000;
    rom[216] = 120'h0D81407E4800000000000D90DA3;
    rom[217] = 120'h0D9300000000000000000000001;
    rom[218] = 120'h0DA300000000000000000000000;
    rom[219] = 120'h0DB1407F4800000000000DC0DD3;
    rom[220] = 120'h0DC300000000000000000000001;
    rom[221] = 120'h0DDA43D14140000000000DE0DF3;
    rom[222] = 120'h0DE300000000000000000000000;
    rom[223] = 120'h0DF300000000000000000000001;
    rom[224] = 120'h0E01407E4800000000000E10E63;
    rom[225] = 120'h0E114079D800000000000E20E53;
    rom[226] = 120'h0E2041D8EC33900000000E30E43;
    rom[227] = 120'h0E3300000000000000000000000;
    rom[228] = 120'h0E4300000000000000000000000;
    rom[229] = 120'h0E5300000000000000000000001;
    rom[230] = 120'h0E6A43E6F906A00000000E70EA3;
    rom[231] = 120'h0E71407E6800000000000E80E93;
    rom[232] = 120'h0E8300000000000000000000000;
    rom[233] = 120'h0E9300000000000000000000000;
    rom[234] = 120'h0EA300000000000000000000001;
    rom[235] = 120'h0EB140799800000000000EC0F53;
    rom[236] = 120'h0EC041D8EC33800000000ED0F43;
    rom[237] = 120'h0ED041D8EC33500000000EE0F13;
    rom[238] = 120'h0EEA43EBBAF8F00000000EF0F03;
    rom[239] = 120'h0EF300000000000000000000000;
    rom[240] = 120'h0F0300000000000000000000001;
    rom[241] = 120'h0F1A43EC2932B00000000F20F33;
    rom[242] = 120'h0F2300000000000000000000000;
    rom[243] = 120'h0F3300000000000000000000001;
    rom[244] = 120'h0F4300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
