module tree_rom_20 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000140681000000000000010023;
    rom[1] = 120'h001300000000000000000000001;
    rom[2] = 120'h002A43D3FFE4D00000000030C23;
    rom[3] = 120'h003A43600000C000000000405F3;
    rom[4] = 120'h004041D8EC33900000000050403;
    rom[5] = 120'h005041D8EC33500000000060233;
    rom[6] = 120'h006A417007B4E00000000070143;
    rom[7] = 120'h007A41391EFA0000000000800F3;
    rom[8] = 120'h0081406890000000000000900C3;
    rom[9] = 120'h0091406830000000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00C1408A54000000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00F1408A5800000000000100133;
    rom[16] = 120'h0101408A3800000000000110123;
    rom[17] = 120'h011300000000000000000000001;
    rom[18] = 120'h012300000000000000000000000;
    rom[19] = 120'h013300000000000000000000001;
    rom[20] = 120'h0141407E18000000000001501C3;
    rom[21] = 120'h015A41EF885EE00000000160193;
    rom[22] = 120'h0161406E1000000000000170183;
    rom[23] = 120'h017300000000000000000000001;
    rom[24] = 120'h018300000000000000000000000;
    rom[25] = 120'h0191407838000000000001A01B3;
    rom[26] = 120'h01A300000000000000000000000;
    rom[27] = 120'h01B300000000000000000000000;
    rom[28] = 120'h01CA41994880A000000001D0203;
    rom[29] = 120'h01D1408B1C000000000001E01F3;
    rom[30] = 120'h01E300000000000000000000000;
    rom[31] = 120'h01F300000000000000000000001;
    rom[32] = 120'h02014087D000000000000210223;
    rom[33] = 120'h021300000000000000000000001;
    rom[34] = 120'h022300000000000000000000001;
    rom[35] = 120'h0231408A5400000000000240333;
    rom[36] = 120'h024A432257EA2000000002502C3;
    rom[37] = 120'h0251406E1000000000000260293;
    rom[38] = 120'h026041D8EC33700000000270283;
    rom[39] = 120'h027300000000000000000000001;
    rom[40] = 120'h028300000000000000000000001;
    rom[41] = 120'h0291407F38000000000002A02B3;
    rom[42] = 120'h02A300000000000000000000000;
    rom[43] = 120'h02B300000000000000000000000;
    rom[44] = 120'h02C041D8EC337000000002D0303;
    rom[45] = 120'h02DA432400181000000002E02F3;
    rom[46] = 120'h02E300000000000000000000001;
    rom[47] = 120'h02F300000000000000000000001;
    rom[48] = 120'h030140691000000000000310323;
    rom[49] = 120'h031300000000000000000000000;
    rom[50] = 120'h032300000000000000000000001;
    rom[51] = 120'h033A3FE00000000000000340393;
    rom[52] = 120'h03414099A600000000000350383;
    rom[53] = 120'h035041D8EC33700000000360373;
    rom[54] = 120'h036300000000000000000000000;
    rom[55] = 120'h037300000000000000000000000;
    rom[56] = 120'h038300000000000000000000000;
    rom[57] = 120'h039041D8EC337000000003A03D3;
    rom[58] = 120'h03AA426C2450F000000003B03C3;
    rom[59] = 120'h03B300000000000000000000001;
    rom[60] = 120'h03C300000000000000000000001;
    rom[61] = 120'h03D1408FC4000000000003E03F3;
    rom[62] = 120'h03E300000000000000000000001;
    rom[63] = 120'h03F300000000000000000000001;
    rom[64] = 120'h040041D8EC33B00000000410563;
    rom[65] = 120'h0411406BA000000000000420493;
    rom[66] = 120'h042A419C0082100000000430483;
    rom[67] = 120'h043A40C00800000000000440453;
    rom[68] = 120'h044300000000000000000000001;
    rom[69] = 120'h045A418C0104200000000460473;
    rom[70] = 120'h046300000000000000000000000;
    rom[71] = 120'h047300000000000000000000001;
    rom[72] = 120'h048300000000000000000000000;
    rom[73] = 120'h049A41EFF1500000000004A04F3;
    rom[74] = 120'h04A14075F8000000000004B04E3;
    rom[75] = 120'h04BA41943E059200000004C04D3;
    rom[76] = 120'h04C300000000000000000000000;
    rom[77] = 120'h04D300000000000000000000000;
    rom[78] = 120'h04E300000000000000000000000;
    rom[79] = 120'h04FA41F80000000000000500533;
    rom[80] = 120'h05014085B400000000000510523;
    rom[81] = 120'h051300000000000000000000000;
    rom[82] = 120'h052300000000000000000000001;
    rom[83] = 120'h053A42CFC084A00000000540553;
    rom[84] = 120'h054300000000000000000000000;
    rom[85] = 120'h055300000000000000000000000;
    rom[86] = 120'h056A421C0000000000000570583;
    rom[87] = 120'h057300000000000000000000000;
    rom[88] = 120'h058041D8EC33F000000005905E3;
    rom[89] = 120'h059041D8EC33D000000005A05B3;
    rom[90] = 120'h05A300000000000000000000000;
    rom[91] = 120'h05BA422500000000000005C05D3;
    rom[92] = 120'h05C300000000000000000000001;
    rom[93] = 120'h05D300000000000000000000000;
    rom[94] = 120'h05E300000000000000000000000;
    rom[95] = 120'h05FA43A0B44FB000000006008D3;
    rom[96] = 120'h0601408FCC000000000006107C3;
    rom[97] = 120'h061041D8EC337000000006206F3;
    rom[98] = 120'h0621407F68000000000006306A3;
    rom[99] = 120'h06314077C000000000000640673;
    rom[100] = 120'h064A4360815FA00000000650663;
    rom[101] = 120'h065300000000000000000000000;
    rom[102] = 120'h066300000000000000000000000;
    rom[103] = 120'h067A436F0FB4B00000000680693;
    rom[104] = 120'h068300000000000000000000001;
    rom[105] = 120'h069300000000000000000000000;
    rom[106] = 120'h06A1408E04000000000006B06C3;
    rom[107] = 120'h06B300000000000000000000001;
    rom[108] = 120'h06CA4374B0000000000006D06E3;
    rom[109] = 120'h06D300000000000000000000001;
    rom[110] = 120'h06E300000000000000000000000;
    rom[111] = 120'h06F1406E9000000000000700753;
    rom[112] = 120'h070A43600600200000000710723;
    rom[113] = 120'h071300000000000000000000000;
    rom[114] = 120'h07214068C000000000000730743;
    rom[115] = 120'h073300000000000000000000000;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h0751407F6000000000000760793;
    rom[118] = 120'h076041D8EC33900000000770783;
    rom[119] = 120'h077300000000000000000000000;
    rom[120] = 120'h078300000000000000000000000;
    rom[121] = 120'h079A436760BD4000000007A07B3;
    rom[122] = 120'h07A300000000000000000000000;
    rom[123] = 120'h07B300000000000000000000000;
    rom[124] = 120'h07C041D8EC339000000007D08C3;
    rom[125] = 120'h07D041D8EC337000000007E0853;
    rom[126] = 120'h07E041D8EC335000000007F0823;
    rom[127] = 120'h07F14093C800000000000800813;
    rom[128] = 120'h080300000000000000000000001;
    rom[129] = 120'h081300000000000000000000001;
    rom[130] = 120'h08214093C600000000000830843;
    rom[131] = 120'h083300000000000000000000001;
    rom[132] = 120'h084300000000000000000000001;
    rom[133] = 120'h085A437B08DE700000000860893;
    rom[134] = 120'h086A4368173CD00000000870883;
    rom[135] = 120'h087300000000000000000000001;
    rom[136] = 120'h088300000000000000000000001;
    rom[137] = 120'h089A437D18F3B000000008A08B3;
    rom[138] = 120'h08A300000000000000000000000;
    rom[139] = 120'h08B300000000000000000000001;
    rom[140] = 120'h08C300000000000000000000000;
    rom[141] = 120'h08D1407E98000000000008E0AB3;
    rom[142] = 120'h08E14068B0000000000008F09C3;
    rom[143] = 120'h08F041D8EC33500000000900973;
    rom[144] = 120'h090A43CA7D45B00000000910943;
    rom[145] = 120'h091140683000000000000920933;
    rom[146] = 120'h092300000000000000000000000;
    rom[147] = 120'h093300000000000000000000000;
    rom[148] = 120'h094A43CC770D500000000950963;
    rom[149] = 120'h095300000000000000000000001;
    rom[150] = 120'h096300000000000000000000001;
    rom[151] = 120'h097041D8EC339000000009809B3;
    rom[152] = 120'h098A43D0162B4000000009909A3;
    rom[153] = 120'h099300000000000000000000000;
    rom[154] = 120'h09A300000000000000000000001;
    rom[155] = 120'h09B300000000000000000000000;
    rom[156] = 120'h09CA43CFF997D000000009D0A43;
    rom[157] = 120'h09D1407988000000000009E0A13;
    rom[158] = 120'h09E1407908000000000009F0A03;
    rom[159] = 120'h09F300000000000000000000001;
    rom[160] = 120'h0A0300000000000000000000001;
    rom[161] = 120'h0A1A43B1D2A2300000000A20A33;
    rom[162] = 120'h0A2300000000000000000000000;
    rom[163] = 120'h0A3300000000000000000000001;
    rom[164] = 120'h0A4A43D17E79E00000000A50A83;
    rom[165] = 120'h0A5A43D01818900000000A60A73;
    rom[166] = 120'h0A6300000000000000000000000;
    rom[167] = 120'h0A7300000000000000000000001;
    rom[168] = 120'h0A8041D8EC33700000000A90AA3;
    rom[169] = 120'h0A9300000000000000000000000;
    rom[170] = 120'h0AA300000000000000000000000;
    rom[171] = 120'h0ABA43D007FE700000000AC0B93;
    rom[172] = 120'h0AC041D8EC33900000000AD0B43;
    rom[173] = 120'h0ADA43AA94B1200000000AE0B13;
    rom[174] = 120'h0AEA43AA0517E00000000AF0B03;
    rom[175] = 120'h0AF300000000000000000000001;
    rom[176] = 120'h0B0300000000000000000000001;
    rom[177] = 120'h0B11407F5800000000000B20B33;
    rom[178] = 120'h0B2300000000000000000000001;
    rom[179] = 120'h0B3300000000000000000000001;
    rom[180] = 120'h0B4140915400000000000B50B83;
    rom[181] = 120'h0B5140877800000000000B60B73;
    rom[182] = 120'h0B6300000000000000000000000;
    rom[183] = 120'h0B7300000000000000000000000;
    rom[184] = 120'h0B8300000000000000000000000;
    rom[185] = 120'h0B9140945200000000000BA0C13;
    rom[186] = 120'h0BAA43D10531A00000000BB0BE3;
    rom[187] = 120'h0BBA43D0FF78C00000000BC0BD3;
    rom[188] = 120'h0BC300000000000000000000000;
    rom[189] = 120'h0BD300000000000000000000000;
    rom[190] = 120'h0BEA43D1CC3CC00000000BF0C03;
    rom[191] = 120'h0BF300000000000000000000001;
    rom[192] = 120'h0C0300000000000000000000001;
    rom[193] = 120'h0C1300000000000000000000001;
    rom[194] = 120'h0C2041D8EC33900000000C31023;
    rom[195] = 120'h0C3041D8EC33700000000C40E73;
    rom[196] = 120'h0C4A43DEDBB4700000000C50D43;
    rom[197] = 120'h0C5A43D46D85D00000000C60CD3;
    rom[198] = 120'h0C6041D8EC33500000000C70CC3;
    rom[199] = 120'h0C71407A3000000000000C80CB3;
    rom[200] = 120'h0C8140798000000000000C90CA3;
    rom[201] = 120'h0C9300000000000000000000001;
    rom[202] = 120'h0CA300000000000000000000000;
    rom[203] = 120'h0CB300000000000000000000001;
    rom[204] = 120'h0CC300000000000000000000001;
    rom[205] = 120'h0CD140799800000000000CE0D33;
    rom[206] = 120'h0CEA43D5BA5F700000000CF0D03;
    rom[207] = 120'h0CF300000000000000000000001;
    rom[208] = 120'h0D0041D8EC33500000000D10D23;
    rom[209] = 120'h0D1300000000000000000000001;
    rom[210] = 120'h0D2300000000000000000000001;
    rom[211] = 120'h0D3300000000000000000000001;
    rom[212] = 120'h0D41407F1800000000000D50E23;
    rom[213] = 120'h0D5140798800000000000D60DB3;
    rom[214] = 120'h0D6A43DF6784500000000D70DA3;
    rom[215] = 120'h0D7A43DF1C29B00000000D80D93;
    rom[216] = 120'h0D8300000000000000000000000;
    rom[217] = 120'h0D9300000000000000000000000;
    rom[218] = 120'h0DA300000000000000000000001;
    rom[219] = 120'h0DB14079D800000000000DC0DF3;
    rom[220] = 120'h0DCA43EB4F93600000000DD0DE3;
    rom[221] = 120'h0DD300000000000000000000000;
    rom[222] = 120'h0DE300000000000000000000001;
    rom[223] = 120'h0DF041D8EC33500000000E00E13;
    rom[224] = 120'h0E0300000000000000000000001;
    rom[225] = 120'h0E1300000000000000000000001;
    rom[226] = 120'h0E2A43E00011900000000E30E63;
    rom[227] = 120'h0E3A43DFFF3FA00000000E40E53;
    rom[228] = 120'h0E4300000000000000000000001;
    rom[229] = 120'h0E5300000000000000000000000;
    rom[230] = 120'h0E6300000000000000000000001;
    rom[231] = 120'h0E7A43DFFD1AF00000000E80EF3;
    rom[232] = 120'h0E8140799800000000000E90EE3;
    rom[233] = 120'h0E9140797800000000000EA0EB3;
    rom[234] = 120'h0EA300000000000000000000001;
    rom[235] = 120'h0EBA7FF00000000000000EC0ED3;
    rom[236] = 120'h0EC300000000000000000000000;
    rom[237] = 120'h0ED300000000000000000000001;
    rom[238] = 120'h0EE300000000000000000000001;
    rom[239] = 120'h0EFA43E2016FA00000000F00F73;
    rom[240] = 120'h0F0140902600000000000F10F63;
    rom[241] = 120'h0F114078B000000000000F20F33;
    rom[242] = 120'h0F2300000000000000000000001;
    rom[243] = 120'h0F3A43E01C5F100000000F40F53;
    rom[244] = 120'h0F4300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
