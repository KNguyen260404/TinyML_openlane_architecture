module tree_rom_3 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000A43C2154C500000000010B63;
    rom[1] = 120'h0011408E8C000000000000207F3;
    rom[2] = 120'h002041D8EC33900000000030603;
    rom[3] = 120'h003041D8EC33500000000040313;
    rom[4] = 120'h004140689000000000000050183;
    rom[5] = 120'h005A436EC661C000000000600F3;
    rom[6] = 120'h006140681000000000000070083;
    rom[7] = 120'h007300000000000000000000001;
    rom[8] = 120'h008A4203FB67E000000000900C3;
    rom[9] = 120'h0091406830000000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00CA42419DE58000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000000;
    rom[15] = 120'h00F140681000000000000100113;
    rom[16] = 120'h010300000000000000000000001;
    rom[17] = 120'h011A43AC3CED700000000120153;
    rom[18] = 120'h012A43901FCCA80000000130143;
    rom[19] = 120'h013300000000000000000000000;
    rom[20] = 120'h014300000000000000000000001;
    rom[21] = 120'h015A43C0C6E2B00000000160173;
    rom[22] = 120'h016300000000000000000000000;
    rom[23] = 120'h017300000000000000000000000;
    rom[24] = 120'h018A3FE00000000000000190223;
    rom[25] = 120'h0191408C58000000000001A0213;
    rom[26] = 120'h01A1408014000000000001B01E3;
    rom[27] = 120'h01B1407C18000000000001C01D3;
    rom[28] = 120'h01C300000000000000000000000;
    rom[29] = 120'h01D300000000000000000000000;
    rom[30] = 120'h01E14088D8000000000001F0203;
    rom[31] = 120'h01F300000000000000000000001;
    rom[32] = 120'h020300000000000000000000000;
    rom[33] = 120'h021300000000000000000000001;
    rom[34] = 120'h0221407E58000000000002302A3;
    rom[35] = 120'h023A41EF934BC00000000240273;
    rom[36] = 120'h024A41DFC65E000000000250263;
    rom[37] = 120'h025300000000000000000000000;
    rom[38] = 120'h026300000000000000000000001;
    rom[39] = 120'h027A43B384412000000000280293;
    rom[40] = 120'h028300000000000000000000000;
    rom[41] = 120'h029300000000000000000000000;
    rom[42] = 120'h02AA437003D72000000002B02E3;
    rom[43] = 120'h02BA416D501EA000000002C02D3;
    rom[44] = 120'h02C300000000000000000000001;
    rom[45] = 120'h02D300000000000000000000001;
    rom[46] = 120'h02E1407F58000000000002F0303;
    rom[47] = 120'h02F300000000000000000000000;
    rom[48] = 120'h030300000000000000000000001;
    rom[49] = 120'h031041D8EC33700000000320433;
    rom[50] = 120'h032140681000000000000330343;
    rom[51] = 120'h033300000000000000000000001;
    rom[52] = 120'h034A436000A11000000003503C3;
    rom[53] = 120'h0351406E1000000000000360393;
    rom[54] = 120'h03614068B000000000000370383;
    rom[55] = 120'h037300000000000000000000000;
    rom[56] = 120'h038300000000000000000000001;
    rom[57] = 120'h039A431CD5C04000000003A03B3;
    rom[58] = 120'h03A300000000000000000000000;
    rom[59] = 120'h03B300000000000000000000001;
    rom[60] = 120'h03C1407E98000000000003D0403;
    rom[61] = 120'h03D14068B0000000000003E03F3;
    rom[62] = 120'h03E300000000000000000000000;
    rom[63] = 120'h03F300000000000000000000000;
    rom[64] = 120'h0401408E0400000000000410423;
    rom[65] = 120'h041300000000000000000000001;
    rom[66] = 120'h042300000000000000000000000;
    rom[67] = 120'h0431407E1800000000000440533;
    rom[68] = 120'h0441406E10000000000004504C3;
    rom[69] = 120'h045A42F4B75A700000000460493;
    rom[70] = 120'h04614068C000000000000470483;
    rom[71] = 120'h047300000000000000000000001;
    rom[72] = 120'h048300000000000000000000001;
    rom[73] = 120'h0491406800000000000004A04B3;
    rom[74] = 120'h04A300000000000000000000001;
    rom[75] = 120'h04B300000000000000000000000;
    rom[76] = 120'h04CA43B0B07F1000000004D0503;
    rom[77] = 120'h04DA43664BBAA000000004E04F3;
    rom[78] = 120'h04E300000000000000000000000;
    rom[79] = 120'h04F300000000000000000000000;
    rom[80] = 120'h050A43B8AD91900000000510523;
    rom[81] = 120'h051300000000000000000000001;
    rom[82] = 120'h052300000000000000000000001;
    rom[83] = 120'h053A42A27843C00000000540593;
    rom[84] = 120'h0541408A5800000000000550583;
    rom[85] = 120'h055A3FF00000000000000560573;
    rom[86] = 120'h056300000000000000000000000;
    rom[87] = 120'h057300000000000000000000000;
    rom[88] = 120'h058300000000000000000000001;
    rom[89] = 120'h0591408E00000000000005A05D3;
    rom[90] = 120'h05A1407EA8000000000005B05C3;
    rom[91] = 120'h05B300000000000000000000001;
    rom[92] = 120'h05C300000000000000000000001;
    rom[93] = 120'h05DA4370D183F000000005E05F3;
    rom[94] = 120'h05E300000000000000000000001;
    rom[95] = 120'h05F300000000000000000000000;
    rom[96] = 120'h0601406BA0000000000006106A3;
    rom[97] = 120'h061041D8EC33B00000000620693;
    rom[98] = 120'h062A419C0082100000000630683;
    rom[99] = 120'h063A40C00800000000000640653;
    rom[100] = 120'h064300000000000000000000001;
    rom[101] = 120'h065A418C0104200000000660673;
    rom[102] = 120'h066300000000000000000000000;
    rom[103] = 120'h067300000000000000000000001;
    rom[104] = 120'h068300000000000000000000000;
    rom[105] = 120'h069300000000000000000000000;
    rom[106] = 120'h06AA42D000001000000006B0783;
    rom[107] = 120'h06B14075F8000000000006C0733;
    rom[108] = 120'h06CA42C001000000000006D0703;
    rom[109] = 120'h06D14073C0000000000006E06F3;
    rom[110] = 120'h06E300000000000000000000000;
    rom[111] = 120'h06F300000000000000000000001;
    rom[112] = 120'h070041D8EC33B00000000710723;
    rom[113] = 120'h071300000000000000000000001;
    rom[114] = 120'h072300000000000000000000000;
    rom[115] = 120'h0731408A4800000000000740753;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h075A4201C3DD180000000760773;
    rom[118] = 120'h076300000000000000000000000;
    rom[119] = 120'h077300000000000000000000001;
    rom[120] = 120'h078041D8EC33B000000007907E3;
    rom[121] = 120'h079A43A520081000000007A07B3;
    rom[122] = 120'h07A300000000000000000000000;
    rom[123] = 120'h07BA43AB1B000000000007C07D3;
    rom[124] = 120'h07C300000000000000000000001;
    rom[125] = 120'h07D300000000000000000000000;
    rom[126] = 120'h07E300000000000000000000000;
    rom[127] = 120'h07FA3FE000000000000008008B3;
    rom[128] = 120'h0801409D5E000000000008108A3;
    rom[129] = 120'h08114094C200000000000820893;
    rom[130] = 120'h082140900200000000000830843;
    rom[131] = 120'h083300000000000000000000000;
    rom[132] = 120'h084041D8EC33700000000850883;
    rom[133] = 120'h08514093B400000000000860873;
    rom[134] = 120'h086300000000000000000000001;
    rom[135] = 120'h087300000000000000000000000;
    rom[136] = 120'h088300000000000000000000000;
    rom[137] = 120'h089300000000000000000000001;
    rom[138] = 120'h08A300000000000000000000000;
    rom[139] = 120'h08B14093C6000000000008C0AB3;
    rom[140] = 120'h08C041D8EC33B000000008D0A03;
    rom[141] = 120'h08D041D8EC339000000008E09B3;
    rom[142] = 120'h08E14093C2000000000008F01203;
    rom[143] = 120'h08FA426C19A9000000000900933;
    rom[144] = 120'h0901408FC400000000000910923;
    rom[145] = 120'h091300000000000000000000001;
    rom[146] = 120'h092300000000000000000000001;
    rom[147] = 120'h093041D8EC33700000000940953;
    rom[148] = 120'h094300000000000000000000001;
    rom[149] = 120'h095300000000000000000000001;
    rom[150] = 120'h0120A43747C29000000000970983;
    rom[151] = 120'h097300000000000000000000001;
    rom[152] = 120'h098A43A6D832D400000009909A3;
    rom[153] = 120'h099300000000000000000000000;
    rom[154] = 120'h09A300000000000000000000001;
    rom[155] = 120'h09B1408F68000000000009C09F3;
    rom[156] = 120'h09CA426510004000000009D09E3;
    rom[157] = 120'h09D300000000000000000000001;
    rom[158] = 120'h09E300000000000000000000000;
    rom[159] = 120'h09F300000000000000000000000;
    rom[160] = 120'h0A0041D8EC33D00000000A10A43;
    rom[161] = 120'h0A1A43BBF184C00000000A20A33;
    rom[162] = 120'h0A2300000000000000000000000;
    rom[163] = 120'h0A3300000000000000000000001;
    rom[164] = 120'h0A41408F6800000000000A50AA3;
    rom[165] = 120'h0A5041D8EC33F00000000A60A93;
    rom[166] = 120'h0A6A42A22800000000000A70A83;
    rom[167] = 120'h0A7300000000000000000000001;
    rom[168] = 120'h0A8300000000000000000000000;
    rom[169] = 120'h0A9300000000000000000000000;
    rom[170] = 120'h0AA300000000000000000000000;
    rom[171] = 120'h0ABA43C20FEBF00000000AC0B53;
    rom[172] = 120'h0AC1409DC200000000000AD0AE3;
    rom[173] = 120'h0AD300000000000000000000001;
    rom[174] = 120'h0AE041D8EC33900000000AF0B43;
    rom[175] = 120'h0AF1409DCE00000000000B00B33;
    rom[176] = 120'h0B0A42AFBBE0300000000B10B23;
    rom[177] = 120'h0B1300000000000000000000001;
    rom[178] = 120'h0B2300000000000000000000000;
    rom[179] = 120'h0B3300000000000000000000001;
    rom[180] = 120'h0B4300000000000000000000000;
    rom[181] = 120'h0B5300000000000000000000000;
    rom[182] = 120'h0B6A43C7FFB4800000000B70B83;
    rom[183] = 120'h0B7300000000000000000000001;
    rom[184] = 120'h0B8A43D3FFE4D00000000B90FA3;
    rom[185] = 120'h0B9A43D1B9C1000000000BA0E13;
    rom[186] = 120'h0BA041D8EC33700000000BB0D43;
    rom[187] = 120'h0BBA43C9F29A400000000BC0C53;
    rom[188] = 120'h0BCA43C80068E00000000BD0BE3;
    rom[189] = 120'h0BD300000000000000000000000;
    rom[190] = 120'h0BE041D8EC33500000000BF0C23;
    rom[191] = 120'h0BFA43C83AA8500000000C00C13;
    rom[192] = 120'h0C0300000000000000000000000;
    rom[193] = 120'h0C1300000000000000000000000;
    rom[194] = 120'h0C2A43C898E1300000000C30C43;
    rom[195] = 120'h0C3300000000000000000000000;
    rom[196] = 120'h0C4300000000000000000000000;
    rom[197] = 120'h0C5A43CFFF90900000000C60CD3;
    rom[198] = 120'h0C6A43CA0048B00000000C70CA3;
    rom[199] = 120'h0C71406B1000000000000C80C93;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C9300000000000000000000001;
    rom[202] = 120'h0CA140683000000000000CB0CC3;
    rom[203] = 120'h0CB300000000000000000000001;
    rom[204] = 120'h0CC300000000000000000000001;
    rom[205] = 120'h0CD1407EA800000000000CE0D13;
    rom[206] = 120'h0CEA43D18ABB800000000CF0D03;
    rom[207] = 120'h0CF300000000000000000000000;
    rom[208] = 120'h0D0300000000000000000000001;
    rom[209] = 120'h0D1140932200000000000D20D33;
    rom[210] = 120'h0D2300000000000000000000001;
    rom[211] = 120'h0D3300000000000000000000001;
    rom[212] = 120'h0D4041D8EC33900000000D50E03;
    rom[213] = 120'h0D51407FB800000000000D60DB3;
    rom[214] = 120'h0D614067E000000000000D70D83;
    rom[215] = 120'h0D7300000000000000000000001;
    rom[216] = 120'h0D8A43CA00A7900000000D90DA3;
    rom[217] = 120'h0D9300000000000000000000000;
    rom[218] = 120'h0DA300000000000000000000000;
    rom[219] = 120'h0DBA43D00864100000000DC0DD3;
    rom[220] = 120'h0DC300000000000000000000001;
    rom[221] = 120'h0DDA43D08EBEA00000000DE0DF3;
    rom[222] = 120'h0DE300000000000000000000000;
    rom[223] = 120'h0DF300000000000000000000001;
    rom[224] = 120'h0E0300000000000000000000000;
    rom[225] = 120'h0E11407EA000000000000E20EF3;
    rom[226] = 120'h0E2140729000000000000E30E43;
    rom[227] = 120'h0E3300000000000000000000001;
    rom[228] = 120'h0E4041D8EC33700000000E50EA3;
    rom[229] = 120'h0E5A43D1C13D300000000E60E73;
    rom[230] = 120'h0E6300000000000000000000000;
    rom[231] = 120'h0E7A43D3F183D00000000E80E93;
    rom[232] = 120'h0E8300000000000000000000001;
    rom[233] = 120'h0E9300000000000000000000000;
    rom[234] = 120'h0EA041D8EC33900000000EB0EE3;
    rom[235] = 120'h0EBA43D1CAC2B00000000EC0ED3;
    rom[236] = 120'h0EC300000000000000000000000;
    rom[237] = 120'h0ED300000000000000000000000;
    rom[238] = 120'h0EE300000000000000000000000;
    rom[239] = 120'h0EF041D8EC33900000000F00F93;
    rom[240] = 120'h0F0140944E00000000000F10F23;
    rom[241] = 120'h0F1300000000000000000000001;
    rom[242] = 120'h0F2041D8EC33700000000F30F63;
    rom[243] = 120'h0F3140945200000000000F40F53;
    rom[244] = 120'h0F4300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 

