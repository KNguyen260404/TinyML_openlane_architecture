module tree_rom_8 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000A43C2154C500000000010CC3;
    rom[1] = 120'h0011408E8C00000000000020753;
    rom[2] = 120'h002041D8EC339000000000305A3;
    rom[3] = 120'h003041D8EC33500000000040293;
    rom[4] = 120'h004140689000000000000050103;
    rom[5] = 120'h005140681000000000000060073;
    rom[6] = 120'h006300000000000000000000001;
    rom[7] = 120'h0071406830000000000000800F3;
    rom[8] = 120'h008A4203FB67E000000000900C3;
    rom[9] = 120'h009A403700000000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00CA437505770000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000000;
    rom[15] = 120'h00F300000000000000000000001;
    rom[16] = 120'h010A3FE000000000000001101A3;
    rom[17] = 120'h0111408C5800000000000120193;
    rom[18] = 120'h012140726000000000000130163;
    rom[19] = 120'h013140692000000000000140153;
    rom[20] = 120'h014300000000000000000000000;
    rom[21] = 120'h015300000000000000000000001;
    rom[22] = 120'h016140801400000000000170183;
    rom[23] = 120'h017300000000000000000000000;
    rom[24] = 120'h018300000000000000000000000;
    rom[25] = 120'h019300000000000000000000001;
    rom[26] = 120'h01AA435FFC444000000001B0223;
    rom[27] = 120'h01B1407E18000000000001C01F3;
    rom[28] = 120'h01C1406E10000000000001D01E3;
    rom[29] = 120'h01D300000000000000000000001;
    rom[30] = 120'h01E300000000000000000000000;
    rom[31] = 120'h01FA416FBF5BF00000000200213;
    rom[32] = 120'h020300000000000000000000001;
    rom[33] = 120'h021300000000000000000000001;
    rom[34] = 120'h022A43B1D47E500000000230263;
    rom[35] = 120'h0231407F6800000000000240253;
    rom[36] = 120'h024300000000000000000000000;
    rom[37] = 120'h025300000000000000000000001;
    rom[38] = 120'h02614068B000000000000270283;
    rom[39] = 120'h027300000000000000000000000;
    rom[40] = 120'h028300000000000000000000001;
    rom[41] = 120'h0291407E58000000000002A03B3;
    rom[42] = 120'h02A1406810000000000002B02C3;
    rom[43] = 120'h02B300000000000000000000001;
    rom[44] = 120'h02CA40EFEF900000000002D0343;
    rom[45] = 120'h02D1407338000000000002E0313;
    rom[46] = 120'h02EA40CEAA000000000002F0303;
    rom[47] = 120'h02F300000000000000000000001;
    rom[48] = 120'h030300000000000000000000001;
    rom[49] = 120'h031041D8EC33700000000320333;
    rom[50] = 120'h032300000000000000000000000;
    rom[51] = 120'h033300000000000000000000000;
    rom[52] = 120'h03414077C800000000000350383;
    rom[53] = 120'h035A4360009C400000000360373;
    rom[54] = 120'h036300000000000000000000000;
    rom[55] = 120'h037300000000000000000000000;
    rom[56] = 120'h038041D8EC337000000003903A3;
    rom[57] = 120'h039300000000000000000000000;
    rom[58] = 120'h03A300000000000000000000000;
    rom[59] = 120'h03B041D8EC337000000003C04B3;
    rom[60] = 120'h03C1408614000000000003D0443;
    rom[61] = 120'h03DA3FF000000000000003E0413;
    rom[62] = 120'h03E1408104000000000003F0403;
    rom[63] = 120'h03F300000000000000000000000;
    rom[64] = 120'h040300000000000000000000001;
    rom[65] = 120'h041A43240018100000000420433;
    rom[66] = 120'h042300000000000000000000001;
    rom[67] = 120'h043300000000000000000000001;
    rom[68] = 120'h0441408A5400000000000450483;
    rom[69] = 120'h045A42A495F1D00000000460473;
    rom[70] = 120'h046300000000000000000000000;
    rom[71] = 120'h047300000000000000000000001;
    rom[72] = 120'h048A4374B0000000000004904A3;
    rom[73] = 120'h049300000000000000000000001;
    rom[74] = 120'h04A300000000000000000000000;
    rom[75] = 120'h04B1408614000000000004C0533;
    rom[76] = 120'h04C1407F38000000000004D0503;
    rom[77] = 120'h04D1407F28000000000004E04F3;
    rom[78] = 120'h04E300000000000000000000001;
    rom[79] = 120'h04F300000000000000000000000;
    rom[80] = 120'h0501407F5800000000000510523;
    rom[81] = 120'h051300000000000000000000001;
    rom[82] = 120'h052300000000000000000000001;
    rom[83] = 120'h0531408A5C00000000000540573;
    rom[84] = 120'h054A42B1BBD8800000000550563;
    rom[85] = 120'h055300000000000000000000000;
    rom[86] = 120'h056300000000000000000000001;
    rom[87] = 120'h0571408E0000000000000580593;
    rom[88] = 120'h058300000000000000000000001;
    rom[89] = 120'h059300000000000000000000000;
    rom[90] = 120'h05A041D8EC33B000000005B0743;
    rom[91] = 120'h05B1406BA0000000000005C0633;
    rom[92] = 120'h05CA419C00821000000005D0623;
    rom[93] = 120'h05DA40C008000000000005E05F3;
    rom[94] = 120'h05E300000000000000000000001;
    rom[95] = 120'h05FA418C0104200000000600613;
    rom[96] = 120'h060300000000000000000000000;
    rom[97] = 120'h061300000000000000000000001;
    rom[98] = 120'h062300000000000000000000000;
    rom[99] = 120'h063A42D000002000000006406D3;
    rom[100] = 120'h064A42C400000000000006506C3;
    rom[101] = 120'h0651408A4800000000000660693;
    rom[102] = 120'h066A41301B0F800000000670683;
    rom[103] = 120'h067300000000000000000000000;
    rom[104] = 120'h068300000000000000000000000;
    rom[105] = 120'h069A4201C1B515C0000006A06B3;
    rom[106] = 120'h06A300000000000000000000000;
    rom[107] = 120'h06B300000000000000000000001;
    rom[108] = 120'h06C300000000000000000000001;
    rom[109] = 120'h06D1407EF0000000000006E06F3;
    rom[110] = 120'h06E300000000000000000000000;
    rom[111] = 120'h06F14086D800000000000700733;
    rom[112] = 120'h070A43A13000080000000710723;
    rom[113] = 120'h071300000000000000000000000;
    rom[114] = 120'h072300000000000000000000000;
    rom[115] = 120'h073300000000000000000000000;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h07514094AA00000000000760BD3;
    rom[118] = 120'h076A426C2450F00000000770983;
    rom[119] = 120'h0771408FC400000000000780893;
    rom[120] = 120'h078041D8EC33500000000790803;
    rom[121] = 120'h079A401800000000000007A07B3;
    rom[122] = 120'h07A300000000000000000000000;
    rom[123] = 120'h07B1408F44000000000007C07D3;
    rom[124] = 120'h07C300000000000000000000001;
    rom[125] = 120'h07DA423A6287BF00000007E07F3;
    rom[126] = 120'h07E300000000000000000000001;
    rom[127] = 120'h07F300000000000000000000001;
    rom[128] = 120'h080041D8EC33C00000000810863;
    rom[129] = 120'h0811408F4400000000000820833;
    rom[130] = 120'h082300000000000000000000001;
    rom[131] = 120'h083A40290000000000000840853;
    rom[132] = 120'h084300000000000000000000000;
    rom[133] = 120'h085300000000000000000000001;
    rom[134] = 120'h086A42140000000000000870883;
    rom[135] = 120'h087300000000000000000000000;
    rom[136] = 120'h088300000000000000000000001;
    rom[137] = 120'h089041D8EC339000000008A0973;
    rom[138] = 120'h08AA3FE000000000000008B0903;
    rom[139] = 120'h08B041D8EC337000000008C08F3;
    rom[140] = 120'h08C1409002000000000008D08E3;
    rom[141] = 120'h08D300000000000000000000000;
    rom[142] = 120'h08E300000000000000000000000;
    rom[143] = 120'h08F300000000000000000000000;
    rom[144] = 120'h090A408A4400000000000910943;
    rom[145] = 120'h091041D8EC33700000000920933;
    rom[146] = 120'h092300000000000000000000001;
    rom[147] = 120'h093300000000000000000000000;
    rom[148] = 120'h0941408FCC00000000000950963;
    rom[149] = 120'h095300000000000000000000000;
    rom[150] = 120'h096300000000000000000000001;
    rom[151] = 120'h097300000000000000000000000;
    rom[152] = 120'h098041D8EC33900000000990B43;
    rom[153] = 120'h099041D8EC337000000009A0A73;
    rom[154] = 120'h09A1408FCC000000000009B0A23;
    rom[155] = 120'h09B041D8EC335000000009C09F3;
    rom[156] = 120'h09CA43A96E58D000000009D09E3;
    rom[157] = 120'h09D300000000000000000000000;
    rom[158] = 120'h09E300000000000000000000001;
    rom[159] = 120'h09F1408F4400000000000A00A13;
    rom[160] = 120'h0A0300000000000000000000001;
    rom[161] = 120'h0A1300000000000000000000000;
    rom[162] = 120'h0A2140930200000000000A30A43;
    rom[163] = 120'h0A3300000000000000000000001;
    rom[164] = 120'h0A4140930600000000000A50A63;
    rom[165] = 120'h0A5300000000000000000000000;
    rom[166] = 120'h0A6300000000000000000000001;
    rom[167] = 120'h0A71408F8000000000000A80AD3;
    rom[168] = 120'h0A81408F4000000000000A90AA3;
    rom[169] = 120'h0A9300000000000000000000001;
    rom[170] = 120'h0AAA43B33A1C400000000AB0AC3;
    rom[171] = 120'h0AB300000000000000000000000;
    rom[172] = 120'h0AC300000000000000000000001;
    rom[173] = 120'h0ADA43375153F00000000AE0B13;
    rom[174] = 120'h0AE140933A00000000000AF0B03;
    rom[175] = 120'h0AF300000000000000000000001;
    rom[176] = 120'h0B0300000000000000000000000;
    rom[177] = 120'h0B11408FD400000000000B20B33;
    rom[178] = 120'h0B2300000000000000000000000;
    rom[179] = 120'h0B3300000000000000000000000;
    rom[180] = 120'h0B4041D8EC33D00000000B50BC3;
    rom[181] = 120'h0B5041D8EC33B00000000B60B73;
    rom[182] = 120'h0B6300000000000000000000000;
    rom[183] = 120'h0B71408F6800000000000B80BB3;
    rom[184] = 120'h0B8A43BBF184C00000000B90BA3;
    rom[185] = 120'h0B9300000000000000000000000;
    rom[186] = 120'h0BA300000000000000000000001;
    rom[187] = 120'h0BB300000000000000000000000;
    rom[188] = 120'h0BC300000000000000000000000;
    rom[189] = 120'h0BD1409DC200000000000BE0BF3;
    rom[190] = 120'h0BE300000000000000000000001;
    rom[191] = 120'h0BFA3FE00000000000000C00C13;
    rom[192] = 120'h0C0300000000000000000000000;
    rom[193] = 120'h0C1041D8EC33900000000C20CB3;
    rom[194] = 120'h0C21409DCE00000000000C30CA3;
    rom[195] = 120'h0C3041D8EC33700000000C40C73;
    rom[196] = 120'h0C4041D8EC33500000000C50C63;
    rom[197] = 120'h0C5300000000000000000000000;
    rom[198] = 120'h0C6300000000000000000000000;
    rom[199] = 120'h0C7A4340C111600000000C80C93;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C9300000000000000000000001;
    rom[202] = 120'h0CA300000000000000000000001;
    rom[203] = 120'h0CB300000000000000000000000;
    rom[204] = 120'h0CCA43C7FFA6C00000000CD0CE3;
    rom[205] = 120'h0CD300000000000000000000001;
    rom[206] = 120'h0CEA43D3FFE4D00000000CF0F43;
    rom[207] = 120'h0CF1407F5800000000000D00E93;
    rom[208] = 120'h0D0140681000000000000D10D23;
    rom[209] = 120'h0D1300000000000000000000001;
    rom[210] = 120'h0D21407E9800000000000D30E23;
    rom[211] = 120'h0D3140798800000000000D40DB3;
    rom[212] = 120'h0D414068B000000000000D50D83;
    rom[213] = 120'h0D5041D8EC33500000000D60D73;
    rom[214] = 120'h0D6300000000000000000000000;
    rom[215] = 120'h0D7300000000000000000000000;
    rom[216] = 120'h0D8A43D1B9C9F00000000D90DA3;
    rom[217] = 120'h0D9300000000000000000000001;
    rom[218] = 120'h0DA300000000000000000000000;
    rom[219] = 120'h0DB041D8EC33700000000DC0DF3;
    rom[220] = 120'h0DCA43CFF997D00000000DD0DE3;
    rom[221] = 120'h0DD300000000000000000000001;
    rom[222] = 120'h0DE300000000000000000000000;
    rom[223] = 120'h0DF041D8EC33900000000E00E13;
    rom[224] = 120'h0E0300000000000000000000000;
    rom[225] = 120'h0E1300000000000000000000000;
    rom[226] = 120'h0E2A43D1380B000000000E30E83;
    rom[227] = 120'h0E31407F4800000000000E40E53;
    rom[228] = 120'h0E4300000000000000000000001;
    rom[229] = 120'h0E5041D8EC33700000000E60E73;
    rom[230] = 120'h0E6300000000000000000000000;
    rom[231] = 120'h0E7300000000000000000000000;
    rom[232] = 120'h0E8300000000000000000000001;
    rom[233] = 120'h0E9041D8EC33900000000EA0F33;
    rom[234] = 120'h0EAA43D0079C500000000EB0EC3;
    rom[235] = 120'h0EB300000000000000000000001;
    rom[236] = 120'h0EC140932200000000000ED0EE3;
    rom[237] = 120'h0ED300000000000000000000001;
    rom[238] = 120'h0EE140945200000000000EF0F23;
    rom[239] = 120'h0EF140932600000000000F00F13;
    rom[240] = 120'h0F0300000000000000000000000;
    rom[241] = 120'h0F1300000000000000000000000;
    rom[242] = 120'h0F2300000000000000000000001;
    rom[243] = 120'h0F3300000000000000000000000;
    rom[244] = 120'h0F4041D8EC33900000000F511E3;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
