module tree_rom_17 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000041D8EC33900000000010BA3;
    rom[1] = 120'h001140681000000000000020033;
    rom[2] = 120'h002300000000000000000000001;
    rom[3] = 120'h0031407F3800000000000040693;
    rom[4] = 120'h004041D8EC335000000000502C3;
    rom[5] = 120'h005A406FD000000000000060133;
    rom[6] = 120'h006A40504000000000000070123;
    rom[7] = 120'h0071406870000000000000800B3;
    rom[8] = 120'h008A403700000000000000900A3;
    rom[9] = 120'h009300000000000000000000001;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B14077E0000000000000C00F3;
    rom[12] = 120'h00CA400800000000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00FA3FF80000000000000100113;
    rom[16] = 120'h010300000000000000000000000;
    rom[17] = 120'h011300000000000000000000001;
    rom[18] = 120'h012300000000000000000000001;
    rom[19] = 120'h0131406930000000000001401D3;
    rom[20] = 120'h014A43CC0B3A5000000001501C3;
    rom[21] = 120'h015140683000000000000160193;
    rom[22] = 120'h016A42000002A02C00000170183;
    rom[23] = 120'h017300000000000000000000001;
    rom[24] = 120'h018300000000000000000000000;
    rom[25] = 120'h0191406890000000000001A01B3;
    rom[26] = 120'h01A300000000000000000000001;
    rom[27] = 120'h01B300000000000000000000000;
    rom[28] = 120'h01C300000000000000000000001;
    rom[29] = 120'h01D14077C8000000000001E0253;
    rom[30] = 120'h01E1406F30000000000001F0223;
    rom[31] = 120'h01F1406E1000000000000200213;
    rom[32] = 120'h020300000000000000000000001;
    rom[33] = 120'h021300000000000000000000000;
    rom[34] = 120'h022A40B27A00000000000230243;
    rom[35] = 120'h023300000000000000000000000;
    rom[36] = 120'h024300000000000000000000001;
    rom[37] = 120'h025A43915644080000000260293;
    rom[38] = 120'h026A43230018000000000270283;
    rom[39] = 120'h027300000000000000000000000;
    rom[40] = 120'h028300000000000000000000001;
    rom[41] = 120'h029A43EA3F08A000000002A02B3;
    rom[42] = 120'h02A300000000000000000000000;
    rom[43] = 120'h02B300000000000000000000001;
    rom[44] = 120'h02C041D8EC337000000002D04C3;
    rom[45] = 120'h02DA436000A0A000000002E03D3;
    rom[46] = 120'h02EA43222E403000000002F0363;
    rom[47] = 120'h02FA419AF35E600000000300333;
    rom[48] = 120'h030A40040000000000000310323;
    rom[49] = 120'h031300000000000000000000000;
    rom[50] = 120'h032300000000000000000000001;
    rom[51] = 120'h0331406E1000000000000340353;
    rom[52] = 120'h034300000000000000000000000;
    rom[53] = 120'h035300000000000000000000000;
    rom[54] = 120'h03614068B0000000000003703A3;
    rom[55] = 120'h037140684000000000000380393;
    rom[56] = 120'h038300000000000000000000000;
    rom[57] = 120'h039300000000000000000000000;
    rom[58] = 120'h03A1407E88000000000003B03C3;
    rom[59] = 120'h03B300000000000000000000001;
    rom[60] = 120'h03C300000000000000000000001;
    rom[61] = 120'h03D14068B0000000000003E0453;
    rom[62] = 120'h03E1406830000000000003F0423;
    rom[63] = 120'h03FA43D5F82D500000000400413;
    rom[64] = 120'h040300000000000000000000000;
    rom[65] = 120'h041300000000000000000000001;
    rom[66] = 120'h042140689000000000000430443;
    rom[67] = 120'h043300000000000000000000001;
    rom[68] = 120'h044300000000000000000000000;
    rom[69] = 120'h045140790800000000000460493;
    rom[70] = 120'h046A4396AADEC00000000470483;
    rom[71] = 120'h047300000000000000000000000;
    rom[72] = 120'h048300000000000000000000001;
    rom[73] = 120'h049A43D409749000000004A04B3;
    rom[74] = 120'h04A300000000000000000000000;
    rom[75] = 120'h04B300000000000000000000000;
    rom[76] = 120'h04CA4329C74E0000000004D05A3;
    rom[77] = 120'h04DA43226FD050000000004E0553;
    rom[78] = 120'h04E1406E10000000000004F0523;
    rom[79] = 120'h04FA42F2E9C2D00000000500513;
    rom[80] = 120'h050300000000000000000000001;
    rom[81] = 120'h051300000000000000000000000;
    rom[82] = 120'h052140783800000000000530543;
    rom[83] = 120'h053300000000000000000000000;
    rom[84] = 120'h054300000000000000000000000;
    rom[85] = 120'h055140683000000000000560573;
    rom[86] = 120'h056300000000000000000000000;
    rom[87] = 120'h0571407E7800000000000580593;
    rom[88] = 120'h058300000000000000000000001;
    rom[89] = 120'h059300000000000000000000001;
    rom[90] = 120'h05AA43E20239C000000005B0623;
    rom[91] = 120'h05BA43C1E7384000000005C05F3;
    rom[92] = 120'h05CA436080086000000005D05E3;
    rom[93] = 120'h05D300000000000000000000000;
    rom[94] = 120'h05E300000000000000000000000;
    rom[95] = 120'h05FA43C7BE9F500000000600613;
    rom[96] = 120'h060300000000000000000000001;
    rom[97] = 120'h061300000000000000000000000;
    rom[98] = 120'h062A43E5C192C00000000630663;
    rom[99] = 120'h063140798000000000000640653;
    rom[100] = 120'h064300000000000000000000001;
    rom[101] = 120'h065300000000000000000000001;
    rom[102] = 120'h066A43EA09ED000000000670683;
    rom[103] = 120'h067300000000000000000000000;
    rom[104] = 120'h068300000000000000000000001;
    rom[105] = 120'h069041D8EC337000000006A0933;
    rom[106] = 120'h06AA3FE000000000000006B0783;
    rom[107] = 120'h06B1408930000000000006C06D3;
    rom[108] = 120'h06C300000000000000000000001;
    rom[109] = 120'h06D14090B6000000000006E0733;
    rom[110] = 120'h06E041D8EC335000000006F0723;
    rom[111] = 120'h06F1408C5800000000000700713;
    rom[112] = 120'h070300000000000000000000000;
    rom[113] = 120'h071300000000000000000000000;
    rom[114] = 120'h072300000000000000000000000;
    rom[115] = 120'h07314093B400000000000740753;
    rom[116] = 120'h074300000000000000000000001;
    rom[117] = 120'h075041D8EC33500000000760773;
    rom[118] = 120'h076300000000000000000000000;
    rom[119] = 120'h077300000000000000000000000;
    rom[120] = 120'h078041D8EC33500000000790863;
    rom[121] = 120'h079A43B0C51BB000000007A0813;
    rom[122] = 120'h07AA436FE82AC000000007B07E3;
    rom[123] = 120'h07B1408A54000000000007C07D3;
    rom[124] = 120'h07C300000000000000000000001;
    rom[125] = 120'h07D300000000000000000000001;
    rom[126] = 120'h07EA43763F613000000007F0803;
    rom[127] = 120'h07F300000000000000000000000;
    rom[128] = 120'h080300000000000000000000000;
    rom[129] = 120'h081A43E00094B00000000820853;
    rom[130] = 120'h08214094AA00000000000830843;
    rom[131] = 120'h083300000000000000000000001;
    rom[132] = 120'h084300000000000000000000001;
    rom[133] = 120'h085300000000000000000000001;
    rom[134] = 120'h086A43A2E867E000000008708E3;
    rom[135] = 120'h0871408E8C000000000008808B3;
    rom[136] = 120'h088A41702EE5D800000008908A3;
    rom[137] = 120'h089300000000000000000000001;
    rom[138] = 120'h08A300000000000000000000000;
    rom[139] = 120'h08B1408FDC000000000008C08D3;
    rom[140] = 120'h08C300000000000000000000001;
    rom[141] = 120'h08D300000000000000000000001;
    rom[142] = 120'h08E14094AA000000000008F0923;
    rom[143] = 120'h08F1408F4400000000000900913;
    rom[144] = 120'h090300000000000000000000001;
    rom[145] = 120'h091300000000000000000000001;
    rom[146] = 120'h092300000000000000000000001;
    rom[147] = 120'h0931408614000000000009409F3;
    rom[148] = 120'h0941407F58000000000009509E3;
    rom[149] = 120'h0951407F4800000000000960973;
    rom[150] = 120'h096300000000000000000000001;
    rom[151] = 120'h097A43A130000800000009809B3;
    rom[152] = 120'h098A43601000400883C509909A3;
    rom[153] = 120'h099300000000000000000000001;
    rom[154] = 120'h09A300000000000000000000000;
    rom[155] = 120'h09BA43B911801000000009C09D3;
    rom[156] = 120'h09C300000000000000000000001;
    rom[157] = 120'h09D300000000000000000000000;
    rom[158] = 120'h09E300000000000000000000001;
    rom[159] = 120'h09FA41A8E047D00000000A00AB3;
    rom[160] = 120'h0A01408A6000000000000A10A63;
    rom[161] = 120'h0A1A400C0000000000000A20A33;
    rom[162] = 120'h0A2300000000000000000000000;
    rom[163] = 120'h0A3A4167CB0FA00000000A40A53;
    rom[164] = 120'h0A4300000000000000000000001;
    rom[165] = 120'h0A5300000000000000000000000;
    rom[166] = 120'h0A6A3FE00000000000000A70A83;
    rom[167] = 120'h0A7300000000000000000000000;
    rom[168] = 120'h0A8A40840400000000000A90AA3;
    rom[169] = 120'h0A9300000000000000000000001;
    rom[170] = 120'h0AA300000000000000000000001;
    rom[171] = 120'h0AB1408E8C00000000000AC0B33;
    rom[172] = 120'h0AC14087CC00000000000AD0B03;
    rom[173] = 120'h0AD14087C400000000000AE0AF3;
    rom[174] = 120'h0AE300000000000000000000000;
    rom[175] = 120'h0AF300000000000000000000000;
    rom[176] = 120'h0B01408E0400000000000B10B23;
    rom[177] = 120'h0B1300000000000000000000001;
    rom[178] = 120'h0B2300000000000000000000000;
    rom[179] = 120'h0B31408F6400000000000B40B73;
    rom[180] = 120'h0B4A43B34813B00000000B50B63;
    rom[181] = 120'h0B5300000000000000000000001;
    rom[182] = 120'h0B6300000000000000000000000;
    rom[183] = 120'h0B7A43E0011B900000000B80B93;
    rom[184] = 120'h0B8300000000000000000000001;
    rom[185] = 120'h0B9300000000000000000000001;
    rom[186] = 120'h0BAA42D00000100000000BB0E43;
    rom[187] = 120'h0BB041D8EC33B00000000BC0D73;
    rom[188] = 120'h0BC1406BA000000000000BD0C43;
    rom[189] = 120'h0BDA419C0082100000000BE0C33;
    rom[190] = 120'h0BEA40C00800000000000BF0C03;
    rom[191] = 120'h0BF300000000000000000000001;
    rom[192] = 120'h0C0A418C0104200000000C10C23;
    rom[193] = 120'h0C1300000000000000000000000;
    rom[194] = 120'h0C2300000000000000000000001;
    rom[195] = 120'h0C3300000000000000000000000;
    rom[196] = 120'h0C41408CCC00000000000C50D03;
    rom[197] = 120'h0C514075F800000000000C60CB3;
    rom[198] = 120'h0C6A42C00100000000000C70CA3;
    rom[199] = 120'h0C714073C000000000000C80C93;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C9300000000000000000000001;
    rom[202] = 120'h0CA300000000000000000000001;
    rom[203] = 120'h0CBA420D9010E00000000CC0CD3;
    rom[204] = 120'h0CC300000000000000000000000;
    rom[205] = 120'h0CDA421EC808700000000CE0CF3;
    rom[206] = 120'h0CE300000000000000000000001;
    rom[207] = 120'h0CF300000000000000000000000;
    rom[208] = 120'h0D0A41E00000270000000D10D23;
    rom[209] = 120'h0D1300000000000000000000000;
    rom[210] = 120'h0D2140917400000000000D30D63;
    rom[211] = 120'h0D3A42651000400000000D40D53;
    rom[212] = 120'h0D4300000000000000000000001;
    rom[213] = 120'h0D5300000000000000000000000;
    rom[214] = 120'h0D6300000000000000000000000;
    rom[215] = 120'h0D71408CCC00000000000D80D93;
    rom[216] = 120'h0D8300000000000000000000000;
    rom[217] = 120'h0D9041D8EC33F00000000DA0E33;
    rom[218] = 120'h0DAA4214000004E000000DB0DC3;
    rom[219] = 120'h0DB300000000000000000000000;
    rom[220] = 120'h0DC140917400000000000DD0E23;
    rom[221] = 120'h0DD041D8EC33D00000000DE0DF3;
    rom[222] = 120'h0DE300000000000000000000000;
    rom[223] = 120'h0DFA42A22800000000000E00E13;
    rom[224] = 120'h0E0300000000000000000000001;
    rom[225] = 120'h0E1300000000000000000000000;
    rom[226] = 120'h0E2300000000000000000000000;
    rom[227] = 120'h0E3300000000000000000000000;
    rom[228] = 120'h0E41407F3000000000000E50E63;
    rom[229] = 120'h0E5300000000000000000000000;
    rom[230] = 120'h0E61408F5800000000000E70F43;
    rom[231] = 120'h0E71408EE800000000000E80F13;
    rom[232] = 120'h0E8041D8EC33B00000000E90F03;
    rom[233] = 120'h0E914086D800000000000EA0EF3;
    rom[234] = 120'h0EAA43A13000080000000EB0EC3;
    rom[235] = 120'h0EB300000000000000000000000;
    rom[236] = 120'h0ECA43AB1B00000000000ED0EE3;
    rom[237] = 120'h0ED300000000000000000000001;
    rom[238] = 120'h0EE300000000000000000000000;
    rom[239] = 120'h0EF300000000000000000000000;
    rom[240] = 120'h0F0300000000000000000000000;
    rom[241] = 120'h0F1A43BBF184C00000000F20F33;
    rom[242] = 120'h0F2300000000000000000000000;
    rom[243] = 120'h0F3300000000000000000000001;
    rom[244] = 120'h0F4300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
