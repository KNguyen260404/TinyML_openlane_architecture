* NGSPICE file created from Random_forest_top_ver2.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VPWR VGND VPB VNB
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__bufinv_16 abstract view
.subckt sky130_fd_sc_hd__bufinv_16 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_1 abstract view
.subckt sky130_fd_sc_hd__clkinv_1 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_4 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinvlp_2 abstract view
.subckt sky130_fd_sc_hd__clkinvlp_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

.subckt Random_forest_top_ver2 VGND VPWR arbitration_id[0] arbitration_id[10] arbitration_id[11]
+ arbitration_id[12] arbitration_id[13] arbitration_id[14] arbitration_id[15] arbitration_id[16]
+ arbitration_id[17] arbitration_id[18] arbitration_id[19] arbitration_id[1] arbitration_id[20]
+ arbitration_id[21] arbitration_id[22] arbitration_id[23] arbitration_id[24] arbitration_id[25]
+ arbitration_id[26] arbitration_id[27] arbitration_id[28] arbitration_id[29] arbitration_id[2]
+ arbitration_id[30] arbitration_id[31] arbitration_id[32] arbitration_id[33] arbitration_id[34]
+ arbitration_id[35] arbitration_id[36] arbitration_id[37] arbitration_id[38] arbitration_id[39]
+ arbitration_id[3] arbitration_id[40] arbitration_id[41] arbitration_id[42] arbitration_id[43]
+ arbitration_id[44] arbitration_id[45] arbitration_id[46] arbitration_id[47] arbitration_id[48]
+ arbitration_id[49] arbitration_id[4] arbitration_id[50] arbitration_id[51] arbitration_id[52]
+ arbitration_id[53] arbitration_id[54] arbitration_id[55] arbitration_id[56] arbitration_id[57]
+ arbitration_id[58] arbitration_id[59] arbitration_id[5] arbitration_id[60] arbitration_id[61]
+ arbitration_id[62] arbitration_id[63] arbitration_id[6] arbitration_id[7] arbitration_id[8]
+ arbitration_id[9] clk data_field[0] data_field[10] data_field[11] data_field[12]
+ data_field[13] data_field[14] data_field[15] data_field[16] data_field[17] data_field[18]
+ data_field[19] data_field[1] data_field[20] data_field[21] data_field[22] data_field[23]
+ data_field[24] data_field[25] data_field[26] data_field[27] data_field[28] data_field[29]
+ data_field[2] data_field[30] data_field[31] data_field[32] data_field[33] data_field[34]
+ data_field[35] data_field[36] data_field[37] data_field[38] data_field[39] data_field[3]
+ data_field[40] data_field[41] data_field[42] data_field[43] data_field[44] data_field[45]
+ data_field[46] data_field[47] data_field[48] data_field[49] data_field[4] data_field[50]
+ data_field[51] data_field[52] data_field[53] data_field[54] data_field[55] data_field[56]
+ data_field[57] data_field[58] data_field[59] data_field[5] data_field[60] data_field[61]
+ data_field[62] data_field[63] data_field[6] data_field[7] data_field[8] data_field[9]
+ feature_valid frame_id_out[0] frame_id_out[1] frame_id_out[2] frame_id_out[3] frame_id_out[4]
+ prediction_out prediction_valid ready_for_next rst_n timestamp[0] timestamp[10]
+ timestamp[11] timestamp[12] timestamp[13] timestamp[14] timestamp[15] timestamp[16]
+ timestamp[17] timestamp[18] timestamp[19] timestamp[1] timestamp[20] timestamp[21]
+ timestamp[22] timestamp[23] timestamp[24] timestamp[25] timestamp[26] timestamp[27]
+ timestamp[28] timestamp[29] timestamp[2] timestamp[30] timestamp[31] timestamp[32]
+ timestamp[33] timestamp[34] timestamp[35] timestamp[36] timestamp[37] timestamp[38]
+ timestamp[39] timestamp[3] timestamp[40] timestamp[41] timestamp[42] timestamp[43]
+ timestamp[44] timestamp[45] timestamp[46] timestamp[47] timestamp[48] timestamp[49]
+ timestamp[4] timestamp[50] timestamp[51] timestamp[52] timestamp[53] timestamp[54]
+ timestamp[55] timestamp[56] timestamp[57] timestamp[58] timestamp[59] timestamp[5]
+ timestamp[60] timestamp[61] timestamp[62] timestamp[63] timestamp[6] timestamp[7]
+ timestamp[8] timestamp[9]
X_3155_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5530__S _1020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6914_ clknet_leaf_70_clk _0627_ net38 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.current_node_data\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6743__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6845_ clknet_leaf_86_clk _0565_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3988_ _1466_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6776_ clknet_leaf_5_clk _0510_ net26 VGND VGND VPWR VPWR complete_votes\[0\] sky130_fd_sc_hd__dfrtp_1
X_5727_ tree_instances\[19\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2772_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5658_ _2703_ _2704_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_92_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4609_ tree_instances\[9\].u_tree.frame_id_out\[4\] tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[9\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5589_ tree_instances\[13\].u_tree.frame_id_out\[0\] current_voting_frame\[0\] VGND
+ VGND VPWR VPWR _2639_ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6484__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire18 _2717_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4960_ _2216_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_47_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3911_ _1391_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_4891_ _1650_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[3\] VGND
+ VGND VPWR VPWR _2171_ sky130_fd_sc_hd__xor2_1
X_6630_ clknet_leaf_57_clk _0389_ net37 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3842_ _1326_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__clkbuf_1
X_6561_ clknet_leaf_50_clk _0335_ net35 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
X_3773_ _1145_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5512_ attack_votes\[4\] VGND VGND VPWR VPWR _2573_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6492_ clknet_leaf_1_clk _0275_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5443_ _2530_ tree_instances\[1\].u_tree.u_tree_weight_rom.gen_tree_1.u_tree_rom.node_data\[12\]
+ _2531_ VGND VGND VPWR VPWR _2532_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5374_ _2461_ VGND VGND VPWR VPWR _2476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_442 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4325_ _1768_ _1789_ VGND VGND VPWR VPWR _1792_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_74_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4256_ _1032_ VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__clkbuf_1
X_4187_ _1652_ VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__clkbuf_1
X_3207_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6995__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6924__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6828_ clknet_leaf_40_clk _0549_ net30 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_93_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6759_ clknet_leaf_4_clk _0000_ net26 VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_46_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_16_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_412 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_14 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_110_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5090_ _1138_ VGND VGND VPWR VPWR _2289_ sky130_fd_sc_hd__inv_2
X_4110_ _1584_ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__clkbuf_1
X_4041_ _1229_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_108_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5992_ _2955_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6335__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4943_ _1727_ _2133_ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6613_ clknet_leaf_36_clk _0377_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
X_4874_ _2146_ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__clkbuf_1
X_3825_ tree_instances\[9\].u_tree.prediction_valid _1025_ VGND VGND VPWR VPWR _1314_
+ sky130_fd_sc_hd__and2b_1
X_6544_ clknet_leaf_43_clk _0318_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3756_ _1247_ _1249_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_76_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6475_ clknet_leaf_99_clk _0263_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5426_ _2521_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3687_ _0858_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__clkbuf_1
X_5357_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _2459_ sky130_fd_sc_hd__inv_2
X_5288_ _2416_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__clkbuf_1
X_4308_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1775_ sky130_fd_sc_hd__inv_2
X_4239_ _1707_ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_71 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4834__A1 _2125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5011__A1 _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6846__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_29_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_104_Right_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3610_ _1123_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__clkbuf_1
X_4590_ _1969_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3541_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6260_ _3129_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3472_ tree_instances\[8\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__buf_2
X_6191_ _0709_ _3035_ VGND VGND VPWR VPWR _3091_ sky130_fd_sc_hd__and2_1
X_5211_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[8\] VGND VGND VPWR
+ VPWR _2376_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5710__C1 _2679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5142_ _2319_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6679__SET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5073_ _2280_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6516__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4024_ _1500_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5975_ _1322_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[1\] tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ _1319_ _2941_ VGND VGND VPWR VPWR _2942_ sky130_fd_sc_hd__a221o_1
X_4926_ _1726_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[6\] _2192_
+ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_82_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4857_ _2139_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__clkbuf_1
X_3808_ _1296_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6527_ clknet_leaf_59_clk _0020_ net38 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4788_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[2\] VGND VGND VPWR
+ VPWR _2091_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3739_ _0976_ _0987_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6458_ clknet_leaf_25_clk _0033_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5409_ _1488_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[1\] VGND
+ VGND VPWR VPWR _2506_ sky130_fd_sc_hd__nand2_1
Xclkload90 clknet_leaf_53_clk VGND VGND VPWR VPWR clkload90/Y sky130_fd_sc_hd__inv_6
X_6389_ clknet_leaf_88_clk _0030_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[2\].u_tree.tree_state\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5684__A net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_367 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6680__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xload_slew30 tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__buf_12
XANTENNA__5471__A1 _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_105_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5760_ _2659_ tree_instances\[6\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2805_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5691_ _2659_ tree_instances\[9\].u_tree.frame_id_out\[3\] tree_instances\[9\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2736_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4711_ _2026_ _2041_ _2042_ _2045_ VGND VGND VPWR VPWR _2046_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_17_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4642_ _1165_ _1999_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ _1595_ VGND VGND VPWR VPWR _2000_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4573_ _1797_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[2\] _1956_
+ VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6312_ clknet_leaf_29_clk _0121_ net28 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3524_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1046_ sky130_fd_sc_hd__buf_1
XFILLER_0_4_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3455_ _0984_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__clkbuf_1
X_6243_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[4\] _2490_ _3116_
+ VGND VGND VPWR VPWR _3121_ sky130_fd_sc_hd__mux2_1
XANTENNA__6768__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3386_ _0920_ _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__nor2_1
X_6174_ _0932_ _3081_ _0038_ tree_instances\[6\].u_tree.pipeline_valid\[0\] VGND VGND
+ VPWR VPWR _0647_ sky130_fd_sc_hd__o2bb2a_1
X_5125_ tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[4\] _2251_ _0018_ VGND
+ VGND VPWR VPWR _2309_ sky130_fd_sc_hd__mux2_1
XANTENNA__6350__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5056_ _2271_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__clkbuf_1
X_4007_ _1484_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_9_Left_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5214__A1 _2122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5958_ _2929_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4909_ tree_instances\[13\].u_tree.read_enable _2188_ VGND VGND VPWR VPWR _2189_
+ sky130_fd_sc_hd__nand2_2
XFILLER_0_47_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5889_ _1400_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[2\] tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ _1395_ _2888_ VGND VGND VPWR VPWR _2889_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5951__B _2553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6438__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_59_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5679__A _2586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6861__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_186 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3240_ _0782_ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__or2_1
X_3171_ _0724_ _0726_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6930_ clknet_leaf_61_clk _0642_ net38 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6861_ clknet_leaf_76_clk _0581_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6792_ clknet_leaf_50_clk _0004_ net34 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5812_ _2844_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5743_ _2586_ _2782_ _2785_ _2787_ VGND VGND VPWR VPWR _2788_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4955__A0 _1832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5674_ tree_instances\[4\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2719_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6949__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4625_ _1784_ _1936_ VGND VGND VPWR VPWR _1987_ sky130_fd_sc_hd__and2_1
X_4556_ _1749_ _1945_ VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3507_ _1028_ _1029_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__nor2_1
XANTENNA__6531__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4487_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND VGND VPWR
+ VPWR _1909_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3438_ _0733_ tree_instances\[7\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _0969_ sky130_fd_sc_hd__or2_1
X_6226_ _0903_ _3109_ _1808_ tree_instances\[5\].u_tree.ready_for_next VGND VGND VPWR
+ VPWR _0671_ sky130_fd_sc_hd__a22o_1
XTAP_TAPCELL_ROW_90_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3369_ _0721_ _0728_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__nor2_1
X_6157_ tree_instances\[1\].u_tree.tree_state\[0\] tree_instances\[1\].u_tree.pipeline_valid\[0\]
+ VGND VGND VPWR VPWR _3067_ sky130_fd_sc_hd__nand2_1
X_5108_ _2300_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__clkbuf_1
X_6088_ _3023_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6094__S _0034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5039_ _1686_ _2222_ VGND VGND VPWR VPWR _2263_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_0_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6619__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput7 net7 VGND VGND VPWR VPWR prediction_out sky130_fd_sc_hd__buf_8
XFILLER_0_31_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_102_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4410_ tree_instances\[7\].u_tree.frame_id_out\[4\] tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[7\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5390_ _2457_ _2482_ VGND VGND VPWR VPWR _2492_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4341_ _1804_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__inv_2
X_4272_ _1738_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6011_ _2965_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5665__A1 _2709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5665__B2 _2708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3223_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5811__S _0004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3154_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0710_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6808__SET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6913_ clknet_leaf_23_clk _0626_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_101 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6844_ clknet_leaf_86_clk _0564_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[8\] sky130_fd_sc_hd__dfrtp_1
X_3987_ _1465_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_99_Left_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6775_ clknet_leaf_5_clk _0509_ net26 VGND VGND VPWR VPWR attack_votes\[4\] sky130_fd_sc_hd__dfrtp_1
X_5726_ _2767_ _2768_ tree_instances\[15\].u_tree.prediction_valid _2770_ VGND VGND
+ VPWR VPWR _2771_ sky130_fd_sc_hd__or4bb_1
XANTENNA__6783__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_79_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5657_ _2691_ _2699_ _2571_ _0000_ VGND VGND VPWR VPWR _2704_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_92_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4608_ _1978_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5588_ _2602_ tree_instances\[13\].u_tree.frame_id_out\[1\] tree_instances\[13\].u_tree.frame_id_out\[2\]
+ _2599_ _2637_ VGND VGND VPWR VPWR _2638_ sky130_fd_sc_hd__a221o_1
X_4539_ tree_instances\[8\].u_tree.frame_id_out\[4\] tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[8\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1942_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_5_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6209_ tree_instances\[5\].u_tree.tree_state\[1\] _3083_ VGND VGND VPWR VPWR _3100_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4395__A1 _1835_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_11_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6453__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3910_ tree_instances\[15\].u_tree.prediction_valid _1137_ VGND VGND VPWR VPWR _1391_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_58_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4890_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[2\] VGND VGND VPWR
+ VPWR _2170_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3841_ _0862_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__clkbuf_1
X_3772_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_532 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6560_ clknet_leaf_3_clk _0334_ net26 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5511_ attack_votes\[0\] attack_votes\[1\] attack_votes\[2\] VGND VGND VPWR VPWR
+ _2572_ sky130_fd_sc_hd__a21oi_1
X_6491_ clknet_leaf_101_clk _0274_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_5442_ _2517_ VGND VGND VPWR VPWR _2531_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5373_ _0944_ VGND VGND VPWR VPWR _2475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4324_ _1776_ VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_74_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_74_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5638__B2 tree_instances\[16\].u_tree.prediction_out VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_4255_ _1716_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__buf_1
X_4186_ _0957_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__clkbuf_1
X_3206_ tree_instances\[20\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__buf_1
XFILLER_0_96_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6964__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6827_ clknet_leaf_41_clk _0548_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6758_ clknet_leaf_66_clk _0493_ net36 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6689_ clknet_leaf_63_clk _0438_ net35 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5709_ _2749_ _2627_ _2750_ _2753_ VGND VGND VPWR VPWR _2754_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6634__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_148 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_26 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4040_ _1514_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5597__A _2578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5991_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[2\] _1431_ _2899_
+ VGND VGND VPWR VPWR _2955_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4942_ _2207_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6612_ clknet_leaf_36_clk _0376_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.prediction_out
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6375__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4873_ _2153_ VGND VGND VPWR VPWR _2154_ sky130_fd_sc_hd__clkbuf_1
X_3824_ _1312_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6304__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6543_ clknet_leaf_42_clk _0317_ net36 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3755_ _1248_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND
+ VPWR VPWR _1249_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_50 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_76_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_289 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6474_ clknet_leaf_9_clk _0262_ net27 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3686_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5425_ _1492_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[1\] _2519_
+ VGND VGND VPWR VPWR _2521_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_12_Right_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5356_ _1248_ VGND VGND VPWR VPWR _2458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5287_ tree_instances\[18\].u_tree.frame_id_out\[1\] tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0753_ VGND VGND VPWR VPWR _2416_ sky130_fd_sc_hd__mux2_1
X_4307_ _1039_ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__buf_1
X_4238_ _1699_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_87_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_94_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_4
X_4169_ _1640_ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_21_Right_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_27_Left_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Right_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_36_Left_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4522__A1 _1837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_85_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_45_Left_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6886__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6815__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4589__A1 _1827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_29_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5538__B1 _1830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_54_Left_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3540_ _1060_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5210_ _2375_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__clkbuf_1
X_3471_ _0731_ tree_instances\[8\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _0999_ sky130_fd_sc_hd__or2_1
X_6190_ _3090_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5710__B1 _2652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5141_ tree_instances\[16\].u_tree.frame_id_out\[4\] tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[16\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2319_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_71_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_63_Left_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5072_ tree_instances\[15\].u_tree.frame_id_out\[4\] tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[15\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2280_ sky130_fd_sc_hd__mux2_1
X_4023_ _0885_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_76_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_92_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6556__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5777__B1 _1020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5974_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[5\] tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ VGND VGND VPWR VPWR _2941_ sky130_fd_sc_hd__xor2_1
XFILLER_0_74_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3252__A1 _0732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4925_ _2198_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_72_Left_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4856_ tree_instances\[12\].u_tree.prediction_out tree_instances\[12\].u_tree.pipeline_prediction\[0\]\[0\]
+ tree_instances\[12\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_30_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3807_ _1295_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6526_ clknet_leaf_59_clk _0019_ net38 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4787_ _2090_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3738_ _0990_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6457_ clknet_leaf_30_clk _0075_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xclkload80 clknet_leaf_44_clk VGND VGND VPWR VPWR clkload80/Y sky130_fd_sc_hd__bufinv_16
X_3669_ _1174_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__clkbuf_1
X_5408_ _0867_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[1\] VGND
+ VGND VPWR VPWR _2505_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_45_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload91 clknet_leaf_54_clk VGND VGND VPWR VPWR clkload91/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6388_ clknet_leaf_86_clk _0029_ net39 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_81_Left_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5339_ complete_votes\[4\] VGND VGND VPWR VPWR _2443_ sky130_fd_sc_hd__inv_2
XANTENNA__6257__A1 _1829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_67_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA__5949__B _2553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_54_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_213 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4743__A1 _1832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_58_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_4
Xload_slew31 tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_12
X_5690_ _2598_ tree_instances\[9\].u_tree.frame_id_out\[0\] tree_instances\[9\].u_tree.frame_id_out\[3\]
+ _2659_ VGND VGND VPWR VPWR _2735_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4710_ _1607_ _1995_ tree_instances\[10\].u_tree.u_tree_weight_rom.cache_valid _2044_
+ _2003_ VGND VGND VPWR VPWR _2045_ sky130_fd_sc_hd__o2111a_1
X_4641_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[4\] VGND VGND VPWR
+ VPWR _1999_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3395__A _0732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4572_ _1959_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6311_ clknet_leaf_29_clk _0120_ net28 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3523_ _1040_ _1044_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3454_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0984_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6242_ _3120_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3385_ _0921_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__clkbuf_1
X_6173_ tree_instances\[6\].u_tree.tree_state\[0\] _0931_ VGND VGND VPWR VPWR _3081_
+ sky130_fd_sc_hd__nand2_1
X_5124_ _2308_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6737__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_49_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_4
X_5055_ tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[1\] _2246_ _0016_ VGND
+ VGND VPWR VPWR _2271_ sky130_fd_sc_hd__mux2_1
X_4006_ _1469_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6390__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_51_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5957_ _1433_ _2553_ VGND VGND VPWR VPWR _2929_ sky130_fd_sc_hd__and2_1
X_4908_ _1686_ _2170_ _2171_ _2187_ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__a211o_1
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5888_ _1409_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[0\] _2885_
+ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR VPWR
+ _2888_ sky130_fd_sc_hd__a2bb2o_1
X_4839_ _2128_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6509_ clknet_leaf_7_clk _0292_ net25 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6478__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6407__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_198 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3170_ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6830__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6860_ clknet_leaf_77_clk _0580_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6791_ clknet_leaf_50_clk _0003_ net35 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5811_ tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[2\] _2595_ _0004_ VGND
+ VGND VPWR VPWR _2844_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5809__S _0004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5742_ _2709_ tree_instances\[14\].u_tree.frame_id_out\[3\] _2786_ tree_instances\[14\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2787_ sky130_fd_sc_hd__o211a_1
XFILLER_0_8_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5673_ _2580_ _2712_ tree_instances\[2\].u_tree.prediction_valid _2715_ net18 VGND
+ VGND VPWR VPWR _2718_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_6_Right_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4624_ _1986_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4555_ _1950_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6989__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3506_ _0843_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6918__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4486_ _1903_ _1904_ _1905_ _1906_ _1907_ VGND VGND VPWR VPWR _1908_ sky130_fd_sc_hd__a221o_1
X_3437_ _0968_ _0965_ tree_instances\[13\].u_tree.tree_state\[1\] VGND VGND VPWR VPWR
+ _0054_ sky130_fd_sc_hd__a21o_1
X_6225_ tree_instances\[5\].u_tree.tree_state\[0\] _0902_ VGND VGND VPWR VPWR _3109_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_90_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _0906_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__clkbuf_1
X_6156_ _2219_ tree_instances\[13\].u_tree.node_data\[12\] _3066_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_data\[12\]
+ _2244_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__a221o_1
X_5107_ _1457_ _2296_ VGND VGND VPWR VPWR _2300_ sky130_fd_sc_hd__and2_1
XANTENNA__6571__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6087_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[6\] _1327_ _3020_
+ VGND VGND VPWR VPWR _3023_ sky130_fd_sc_hd__mux2_1
X_3299_ _0833_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__or2_1
X_5038_ _2262_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_64_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6989_ clknet_leaf_81_clk _0695_ net32 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput8 net8 VGND VGND VPWR VPWR prediction_valid sky130_fd_sc_hd__buf_8
XANTENNA__6659__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5123__A1 _2249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_8_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_102_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_59_Right_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4340_ _1803_ tree_instances\[2\].u_tree.pipeline_valid\[0\] tree_instances\[2\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__or3b_2
XFILLER_0_10_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4271_ _1732_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6329__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6010_ tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[3\] _1834_ _0032_ VGND
+ VGND VPWR VPWR _2965_ sky130_fd_sc_hd__mux2_1
X_3222_ _0771_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__clkbuf_1
X_3153_ _0708_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_68_Right_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_68_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_68_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6912_ clknet_leaf_17_clk _0625_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6843_ clknet_leaf_68_clk _0563_ net39 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3986_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1465_ sky130_fd_sc_hd__inv_2
XPHY_EDGE_ROW_77_Right_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_61_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6774_ clknet_leaf_5_clk _0508_ net26 VGND VGND VPWR VPWR attack_votes\[3\] sky130_fd_sc_hd__dfrtp_1
X_5725_ _2713_ tree_instances\[15\].u_tree.frame_id_out\[1\] tree_instances\[15\].u_tree.frame_id_out\[3\]
+ _2709_ _2769_ VGND VGND VPWR VPWR _2770_ sky130_fd_sc_hd__o221a_1
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5656_ attack_votes\[3\] _2691_ _2699_ VGND VGND VPWR VPWR _2703_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4607_ tree_instances\[9\].u_tree.frame_id_out\[3\] tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _1025_ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_92_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5587_ _2585_ tree_instances\[13\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2637_
+ sky130_fd_sc_hd__xor2_1
X_4538_ _1941_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
X_4469_ _0715_ VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_86_Right_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_5_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6208_ _3099_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6139_ _2104_ _2105_ _2106_ VGND VGND VPWR VPWR _3051_ sky130_fd_sc_hd__nand3_1
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5957__B _2553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_95_Right_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3758__A _0732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_19_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3840_ _1320_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__clkbuf_1
X_3771_ _1260_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5583__B2 _2631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5583__A1 _2579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5510_ attack_votes\[3\] VGND VGND VPWR VPWR _2571_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6490_ clknet_leaf_1_clk _0273_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.cache_valid
+ sky130_fd_sc_hd__dfxtp_1
X_5441_ tree_instances\[1\].u_tree.read_enable VGND VGND VPWR VPWR _2530_ sky130_fd_sc_hd__clkbuf_1
X_5372_ _2463_ VGND VGND VPWR VPWR _2474_ sky130_fd_sc_hd__clkbuf_1
X_4323_ _1777_ VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5638__A2 _2679_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4254_ _1704_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3205_ tree_instances\[2\].u_tree.tree_state\[0\] _0754_ _0755_ VGND VGND VPWR VPWR
+ _0071_ sky130_fd_sc_hd__a21o_1
X_4185_ _1656_ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6826_ clknet_leaf_46_clk _0547_ net36 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.read_enable
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6757_ clknet_leaf_70_clk _0492_ net38 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5708_ tree_instances\[0\].u_tree.frame_id_out\[2\] _2600_ _2751_ _2752_ tree_instances\[0\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2753_ sky130_fd_sc_hd__o221a_1
X_3969_ _1445_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6688_ clknet_leaf_44_clk _0437_ net34 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6933__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5639_ _2653_ _2672_ _2688_ VGND VGND VPWR VPWR _2689_ sky130_fd_sc_hd__nor3_1
XFILLER_0_20_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3463__D tree_instances\[4\].u_tree.ready_for_next VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6674__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6603__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_110_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5990_ _2954_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__clkbuf_1
X_4941_ _1724_ _2133_ VGND VGND VPWR VPWR _2207_ sky130_fd_sc_hd__and2_1
XFILLER_0_24_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4872_ _0810_ VGND VGND VPWR VPWR _2153_ sky130_fd_sc_hd__clkbuf_1
X_6611_ clknet_leaf_36_clk _0375_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3823_ _1311_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6542_ clknet_leaf_45_clk _0316_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3754_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1248_ sky130_fd_sc_hd__buf_1
XFILLER_0_27_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3685_ _1187_ _1189_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_344 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6473_ clknet_leaf_11_clk _0261_ net25 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5424_ _2520_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_76_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_441 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6344__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5355_ _2452_ _0939_ VGND VGND VPWR VPWR _2457_ sky130_fd_sc_hd__nand2_1
X_5286_ _2415_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__clkbuf_1
X_4306_ _1772_ VGND VGND VPWR VPWR _1773_ sky130_fd_sc_hd__clkbuf_1
X_4237_ _1705_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_4_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4168_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1640_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_87_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4099_ _1573_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6809_ clknet_leaf_41_clk _0087_ net36 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_98_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_254 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_100_Left_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5698__A _2588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6855__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_max_cap25_A net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5538__A1 _1827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3470_ _0993_ _0996_ _0998_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__nor3_1
XFILLER_0_51_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5140_ _2318_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5071_ _2279_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__clkbuf_1
X_4022_ _1499_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5973_ _1328_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[3\] tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ _1335_ VGND VGND VPWR VPWR _2940_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_252 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4924_ _1721_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[5\] _2192_
+ VGND VGND VPWR VPWR _2198_ sky130_fd_sc_hd__mux2_1
XANTENNA__6596__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_82_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4855_ _2138_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3806_ _1294_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4786_ _2087_ tree_instances\[12\].u_tree.pipeline_prediction\[0\]\[0\] _2089_ VGND
+ VGND VPWR VPWR _2090_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3737_ _0989_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__clkbuf_1
X_6525_ clknet_leaf_62_clk _0061_ net38 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_43_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload70 clknet_leaf_72_clk VGND VGND VPWR VPWR clkload70/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_15_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3668_ _1173_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__clkbuf_1
X_6456_ clknet_leaf_76_clk _0248_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.gen_tree_20.u_tree_rom.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5407_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND VGND VPWR
+ VPWR _2504_ sky130_fd_sc_hd__inv_2
Xclkload81 clknet_leaf_45_clk VGND VGND VPWR VPWR clkload81/Y sky130_fd_sc_hd__clkinv_2
Xclkload92 clknet_leaf_55_clk VGND VGND VPWR VPWR clkload92/Y sky130_fd_sc_hd__bufinv_16
X_6387_ clknet_leaf_66_clk _0071_ net36 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_11_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3599_ tree_instances\[13\].u_tree.tree_state\[0\] _1113_ _1114_ VGND VGND VPWR VPWR
+ _0053_ sky130_fd_sc_hd__a21o_1
XFILLER_0_100_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5338_ state\[0\] _2441_ VGND VGND VPWR VPWR _2442_ sky130_fd_sc_hd__or2b_1
X_5269_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[6\] _1388_ _2399_
+ VGND VGND VPWR VPWR _2406_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_26_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3469__C tree_instances\[20\].u_tree.ready_for_next VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xload_slew32 tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_12
XANTENNA_clkload6_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5759__A1 _2580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4640_ _1597_ _1995_ _1996_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[7\]
+ _1997_ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6310_ clknet_leaf_29_clk _0119_ net33 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5931__A1 tree_instances\[0\].u_tree.frame_id_in\[4\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_4571_ _1790_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[1\] _1956_
+ VGND VGND VPWR VPWR _1959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3522_ _1043_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3453_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6241_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[3\] _2468_ _3116_
+ VGND VGND VPWR VPWR _3120_ sky130_fd_sc_hd__mux2_1
X_6172_ _3078_ VGND VGND VPWR VPWR _3080_ sky130_fd_sc_hd__clkbuf_1
X_3384_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[3\] tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[2\]
+ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__or2_1
X_5123_ tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[3\] _2249_ _0018_ VGND
+ VGND VPWR VPWR _2308_ sky130_fd_sc_hd__mux2_1
X_5054_ _2270_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4005_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1483_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_84_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6777__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6706__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5956_ _2928_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_23_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_51_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5887_ _1410_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[0\] tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ _1403_ VGND VGND VPWR VPWR _2887_ sky130_fd_sc_hd__a22o_1
X_4907_ _2174_ _2177_ _2181_ _2186_ VGND VGND VPWR VPWR _2187_ sky130_fd_sc_hd__or4_1
XFILLER_0_90_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4838_ tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[4\] _1837_ _0010_ VGND
+ VGND VPWR VPWR _2128_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_556 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4769_ _1615_ _2030_ VGND VGND VPWR VPWR _2080_ sky130_fd_sc_hd__and2_1
XFILLER_0_15_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_95_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6508_ clknet_leaf_1_clk _0291_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_6439_ clknet_leaf_23_clk _0232_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_3_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6447__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_39_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6413__SET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_91_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6790_ clknet_leaf_46_clk _0045_ net34 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XANTENNA_clkbuf_leaf_44_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5810_ _2843_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5741_ _2627_ tree_instances\[14\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2786_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5672_ _2714_ tree_instances\[2\].u_tree.frame_id_out\[2\] tree_instances\[2\].u_tree.frame_id_out\[3\]
+ _2709_ _2716_ VGND VGND VPWR VPWR _2717_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_4_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_59_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4623_ _1764_ _1937_ VGND VGND VPWR VPWR _1986_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4554_ _1759_ _1945_ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_102_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3505_ _1027_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4485_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[7\] tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ VGND VGND VPWR VPWR _1907_ sky130_fd_sc_hd__xor2_1
X_6224_ _3108_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3436_ _0967_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__clkbuf_1
X_3367_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_90_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6155_ _3065_ VGND VGND VPWR VPWR _3066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5106_ _2299_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__clkbuf_1
X_6086_ _3022_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6958__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3298_ _0842_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__clkbuf_1
X_5037_ _1679_ _2222_ VGND VGND VPWR VPWR _2262_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5796__A _2627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6988_ clknet_leaf_95_clk _0694_ net32 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5939_ tree_instances\[2\].u_tree.frame_id_out\[2\] tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0755_ VGND VGND VPWR VPWR _2920_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3466__D tree_instances\[8\].u_tree.ready_for_next VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xoutput9 net22 VGND VGND VPWR VPWR ready_for_next sky130_fd_sc_hd__buf_8
XFILLER_0_9_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6699__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6628__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_3_1__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_48 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4270_ _1737_ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3221_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[5\] tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[4\]
+ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__nor2_1
X_3152_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6369__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_68_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6911_ clknet_leaf_38_clk _0624_ net29 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6842_ clknet_leaf_85_clk _0562_ net39 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3985_ _1463_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_61_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6773_ clknet_leaf_6_clk _0507_ net26 VGND VGND VPWR VPWR attack_votes\[2\] sky130_fd_sc_hd__dfrtp_1
X_5724_ _2603_ tree_instances\[15\].u_tree.frame_id_out\[1\] tree_instances\[15\].u_tree.frame_id_out\[0\]
+ _2598_ VGND VGND VPWR VPWR _2769_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5655_ _1018_ _2701_ _2702_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_79_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4606_ _1977_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5586_ tree_instances\[5\].u_tree.prediction_out _2624_ _2635_ tree_instances\[3\].u_tree.prediction_out
+ VGND VGND VPWR VPWR _2636_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4537_ tree_instances\[8\].u_tree.frame_id_out\[3\] tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _1000_ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4468_ _1890_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3419_ _0951_ _0952_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_5_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6207_ tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[4\] tree_instances\[0\].u_tree.frame_id_in\[4\]
+ _0036_ VGND VGND VPWR VPWR _3099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6792__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4399_ _1838_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_6138_ _2130_ VGND VGND VPWR VPWR _3050_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6721__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6069_ _3009_ VGND VGND VPWR VPWR _3012_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6809__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_19_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3770_ _1144_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5440_ _2528_ VGND VGND VPWR VPWR _2529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5371_ _2472_ VGND VGND VPWR VPWR _2473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4322_ _1773_ _1046_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4253_ _1709_ _1712_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__nor2_1
X_3204_ tree_instances\[2\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__buf_2
X_4184_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1656_ sky130_fd_sc_hd__inv_2
XFILLER_0_96_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6825_ clknet_leaf_39_clk _0546_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6756_ clknet_leaf_24_clk _0491_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3968_ _1054_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__clkbuf_1
X_5707_ tree_instances\[0\].u_tree.frame_id_out\[1\] _2579_ VGND VGND VPWR VPWR _2752_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3899_ _1378_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__clkbuf_1
X_6687_ clknet_leaf_44_clk _0436_ net34 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5638_ tree_instances\[10\].u_tree.prediction_out _2679_ _2687_ tree_instances\[16\].u_tree.prediction_out
+ VGND VGND VPWR VPWR _2688_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5569_ _2599_ VGND VGND VPWR VPWR _2619_ sky130_fd_sc_hd__buf_4
XFILLER_0_103_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6643__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_110_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4940_ _2206_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4871_ _2151_ VGND VGND VPWR VPWR _2152_ sky130_fd_sc_hd__clkbuf_1
X_6610_ clknet_leaf_39_clk _0374_ net30 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3822_ _1006_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6541_ clknet_leaf_1_clk _0315_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.cached_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_54_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3753_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1247_ sky130_fd_sc_hd__inv_2
X_6472_ clknet_leaf_9_clk _0260_ net27 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3684_ _1188_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__buf_1
X_5423_ _1496_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[0\] _2519_
+ VGND VGND VPWR VPWR _2520_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_76_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5354_ _2449_ VGND VGND VPWR VPWR _2456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_453 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4305_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1772_ sky130_fd_sc_hd__inv_2
XFILLER_0_49_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6313__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5285_ tree_instances\[18\].u_tree.frame_id_out\[0\] tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0753_ VGND VGND VPWR VPWR _2415_ sky130_fd_sc_hd__mux2_1
X_4236_ _0839_ _0837_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4167_ _1631_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4098_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1573_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6808_ clknet_leaf_46_clk _0530_ net36 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_41_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6739_ clknet_leaf_70_clk _0487_ net38 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_98_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_49_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6895__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6824__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5338__B_N _2441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5070_ tree_instances\[15\].u_tree.frame_id_out\[3\] tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _1137_ VGND VGND VPWR VPWR _2279_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4021_ tree_instances\[17\].u_tree.prediction_valid _0909_ VGND VGND VPWR VPWR _1499_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5972_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND VGND VPWR
+ VPWR _2939_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4923_ _2197_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_82_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4854_ tree_instances\[12\].u_tree.frame_id_out\[4\] tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[12\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2138_ sky130_fd_sc_hd__mux2_1
X_3805_ _1002_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4785_ _0009_ _2088_ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__or2_1
X_3736_ _0901_ _0894_ _1232_ tree_instances\[19\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0066_ sky130_fd_sc_hd__a31o_1
X_6524_ clknet_leaf_2_clk _0306_ net26 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6565__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6455_ clknet_leaf_24_clk _0089_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
X_3667_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1173_ sky130_fd_sc_hd__buf_1
Xclkload60 clknet_leaf_83_clk VGND VGND VPWR VPWR clkload60/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_30_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload71 clknet_leaf_73_clk VGND VGND VPWR VPWR clkload71/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload82 clknet_leaf_46_clk VGND VGND VPWR VPWR clkload82/Y sky130_fd_sc_hd__bufinv_16
X_6386_ clknet_leaf_55_clk _0192_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload93 clknet_leaf_56_clk VGND VGND VPWR VPWR clkload93/Y sky130_fd_sc_hd__clkinvlp_4
X_5406_ _2503_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__clkbuf_1
X_3598_ tree_instances\[13\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__buf_2
X_5337_ _0731_ _0993_ _0996_ _0998_ VGND VGND VPWR VPWR _2441_ sky130_fd_sc_hd__or4_4
XFILLER_0_11_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5268_ _2405_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4219_ tree_instances\[4\].u_tree.prediction_valid _0849_ VGND VGND VPWR VPWR _1689_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__5799__A _2580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5465__A1 _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5199_ _2328_ _2367_ VGND VGND VPWR VPWR _2370_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_26_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xload_slew33 net36 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__buf_12
XFILLER_0_72_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4570_ _1958_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_515 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3521_ _1041_ _1042_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_25 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_3_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3452_ _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6240_ _3119_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3383_ _0919_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__clkbuf_1
X_6171_ _2561_ VGND VGND VPWR VPWR _3079_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5695__A1 _2576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5695__B2 _2713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_110_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5122_ _2307_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__clkbuf_1
X_5053_ tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[0\] _2122_ _0016_ VGND
+ VGND VPWR VPWR _2270_ sky130_fd_sc_hd__mux2_1
X_4004_ _0871_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_84_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_23_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5955_ _1424_ _2553_ VGND VGND VPWR VPWR _2928_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5886_ _1178_ _2885_ _2882_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[7\]
+ tree_instances\[20\].u_tree.u_tree_weight_rom.cache_valid VGND VGND VPWR VPWR _2886_
+ sky130_fd_sc_hd__o221a_1
X_4906_ _2182_ _2183_ _2184_ _2185_ VGND VGND VPWR VPWR _2186_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4837_ _2127_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4768_ _2079_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3719_ _1216_ _1217_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_95_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6507_ clknet_leaf_1_clk _0290_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_4699_ _2036_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6438_ clknet_leaf_23_clk _0231_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5686__A1 _2713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5686__B2 _2708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6369_ clknet_leaf_19_clk _0176_ net25 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_3_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5041__B _2222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5610__A1 _2659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6487__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5601__A1 _2575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5740_ _2583_ _2783_ tree_instances\[14\].u_tree.frame_id_out\[4\] _2708_ _2784_
+ VGND VGND VPWR VPWR _2785_ sky130_fd_sc_hd__o221a_1
XFILLER_0_57_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6876__CLK clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5671_ _2627_ tree_instances\[2\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2716_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4622_ _1985_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4553_ _1949_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4484_ _1046_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[4\] VGND
+ VGND VPWR VPWR _1906_ sky130_fd_sc_hd__or2_1
X_3504_ _0833_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__clkbuf_1
X_6223_ tree_instances\[5\].u_tree.prediction_out tree_instances\[5\].u_tree.pipeline_prediction\[0\]\[0\]
+ tree_instances\[5\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _3108_ sky130_fd_sc_hd__mux2_1
X_3435_ tree_instances\[13\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__buf_1
XFILLER_0_0_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3366_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_90_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6154_ _3064_ VGND VGND VPWR VPWR _3065_ sky130_fd_sc_hd__clkbuf_1
X_5105_ _1454_ _2296_ VGND VGND VPWR VPWR _2299_ sky130_fd_sc_hd__and2_1
X_6085_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[5\] _1352_ _3020_
+ VGND VGND VPWR VPWR _3022_ sky130_fd_sc_hd__mux2_1
X_3297_ _0836_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__nand2_1
X_5036_ _2261_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6998__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_82 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_69_Left_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_0_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6987_ clknet_leaf_37_clk _0693_ net30 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6927__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5938_ _2919_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3597__A _1112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6580__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5869_ _2875_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_78_Left_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4398__A1 _1837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3220_ _0763_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__nor2_1
X_3151_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_20 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_68_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6910_ clknet_leaf_17_clk _0623_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6841_ clknet_leaf_69_clk _0561_ net39 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6338__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3984_ _1462_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_61_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_33_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6772_ clknet_leaf_5_clk _0506_ net27 VGND VGND VPWR VPWR attack_votes\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5723_ _2576_ tree_instances\[15\].u_tree.frame_id_out\[0\] tree_instances\[15\].u_tree.frame_id_out\[2\]
+ _2714_ VGND VGND VPWR VPWR _2768_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5654_ state\[0\] _2447_ attack_votes\[2\] VGND VGND VPWR VPWR _2702_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_79_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4605_ tree_instances\[9\].u_tree.frame_id_out\[2\] tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _1025_ VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_13_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5585_ _2589_ _2625_ tree_instances\[3\].u_tree.prediction_valid _2626_ _2634_ VGND
+ VGND VPWR VPWR _2635_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4536_ _1940_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4467_ _1889_ VGND VGND VPWR VPWR _1890_ sky130_fd_sc_hd__clkbuf_1
X_3418_ _0733_ tree_instances\[11\].u_tree.pipeline_valid\[0\] tree_instances\[11\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4398_ tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[4\] _1837_ _0040_ VGND
+ VGND VPWR VPWR _1838_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_5_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6206_ _3098_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__clkbuf_1
X_3349_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _0890_ sky130_fd_sc_hd__clkbuf_1
X_6137_ _0909_ _3049_ _0020_ tree_instances\[17\].u_tree.pipeline_valid\[0\] VGND
+ VGND VPWR VPWR _0642_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_84_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5813__A1 _2249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6068_ _3005_ VGND VGND VPWR VPWR _3011_ sky130_fd_sc_hd__clkbuf_1
X_5019_ tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[4\] _2251_ _0014_ VGND
+ VGND VPWR VPWR _2252_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_90_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5600__A _2610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6761__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_527 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_58_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6849__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_619 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_10_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5370_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[8\] VGND VGND VPWR
+ VPWR _2472_ sky130_fd_sc_hd__inv_2
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4543__B2 tree_instances\[8\].u_tree.ready_for_next VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4321_ _1787_ VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__clkbuf_1
X_4252_ _1720_ VGND VGND VPWR VPWR _1721_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_74_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3203_ _0733_ tree_instances\[2\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _0754_ sky130_fd_sc_hd__or2_1
X_4183_ _1650_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6519__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6824_ clknet_leaf_41_clk _0545_ net36 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_6755_ clknet_leaf_25_clk _0050_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3967_ _1062_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5706_ tree_instances\[0\].u_tree.frame_id_out\[1\] _2578_ VGND VGND VPWR VPWR _2751_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_9_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3898_ _1374_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_30_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_4
X_6686_ clknet_leaf_51_clk _0435_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5637_ _2682_ _2683_ _2686_ VGND VGND VPWR VPWR _2687_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5568_ _2600_ tree_instances\[5\].u_tree.frame_id_out\[2\] _2616_ _2617_ tree_instances\[5\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2618_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4519_ _1929_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5499_ _1894_ VGND VGND VPWR VPWR _2564_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_97_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA__6942__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_16_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6100__S _0034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_88_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA__6683__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6612__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_16 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4870_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[8\] VGND VGND VPWR
+ VPWR _2151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3821_ _1292_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6540_ clknet_leaf_4_clk _0314_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_39_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_12_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3752_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[7\] _0945_ VGND VGND
+ VPWR VPWR _1246_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3683_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1188_ sky130_fd_sc_hd__clkbuf_1
X_6471_ clknet_leaf_10_clk _0259_ net25 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5422_ _2518_ VGND VGND VPWR VPWR _2519_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_76_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4516__A1 _1830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5353_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _2455_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6010__S _0032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4304_ _1769_ VGND VGND VPWR VPWR _1771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5284_ _2413_ VGND VGND VPWR VPWR _2414_ sky130_fd_sc_hd__dlymetal6s2s_1
X_4235_ _0840_ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_79_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_4
X_4166_ _1635_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6353__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_87_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4097_ _1567_ VGND VGND VPWR VPWR _1572_ sky130_fd_sc_hd__clkbuf_1
X_6807_ clknet_leaf_45_clk _0529_ net34 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4999_ _2238_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6738_ clknet_leaf_68_clk _0486_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.prediction_out
+ sky130_fd_sc_hd__dfrtp_1
X_6669_ clknet_leaf_63_clk _0419_ net35 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_21_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_98_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5763__A1_N _2600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6962__SET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_14_Left_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_176 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_23_Left_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_552 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6864__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_71_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4020_ _1490_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_1_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_32_Left_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5971_ _1323_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[2\] VGND
+ VGND VPWR VPWR _2938_ sky130_fd_sc_hd__xor2_1
X_4922_ _1727_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[4\] _2192_
+ VGND VGND VPWR VPWR _2197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_82_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4853_ _2137_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3804_ _1003_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__clkbuf_1
X_4784_ tree_instances\[12\].u_tree.tree_state\[0\] tree_instances\[12\].u_tree.tree_state\[1\]
+ tree_instances\[12\].u_tree.tree_state\[2\] _0830_ VGND VGND VPWR VPWR _2088_ sky130_fd_sc_hd__o31ai_1
X_3735_ _1228_ _1231_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6523_ clknet_leaf_7_clk _0091_ net25 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
X_6454_ clknet_leaf_24_clk _0247_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XPHY_EDGE_ROW_41_Left_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload50 clknet_leaf_34_clk VGND VGND VPWR VPWR clkload50/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_70_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3666_ _1172_ _0379_ tree_instances\[10\].u_tree.tree_state\[1\] VGND VGND VPWR VPWR
+ _0048_ sky130_fd_sc_hd__a21o_1
Xclkload61 clknet_leaf_84_clk VGND VGND VPWR VPWR clkload61/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_30_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5405_ tree_instances\[20\].u_tree.u_tree_weight_rom.cache_valid _2502_ VGND VGND
+ VPWR VPWR _2503_ sky130_fd_sc_hd__or2_1
Xclkload83 clknet_leaf_47_clk VGND VGND VPWR VPWR clkload83/Y sky130_fd_sc_hd__inv_6
Xclkload94 clknet_leaf_57_clk VGND VGND VPWR VPWR clkload94/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6385_ clknet_leaf_13_clk _0107_ net29 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3597_ _1112_ tree_instances\[13\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _1113_ sky130_fd_sc_hd__or2_1
Xclkload72 clknet_leaf_74_clk VGND VGND VPWR VPWR clkload72/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5336_ _1252_ _1989_ _1825_ tree_instances\[19\].u_tree.ready_for_next VGND VGND
+ VPWR VPWR _0449_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5267_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[5\] _1383_ _2399_
+ VGND VGND VPWR VPWR _2405_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4218_ _1688_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5799__B _2583_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5198_ _2369_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__clkbuf_1
X_4149_ _1117_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_50_Left_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_26_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_54_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_54_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5039__B _2222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload0 clknet_3_0__leaf_clk VGND VGND VPWR VPWR clkload0/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6796__D _0010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_load_slew37_A net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xload_slew34 net35 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__buf_12
XFILLER_0_96_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_235 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3520_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3451_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _0981_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3382_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[1\] tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[0\]
+ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__or2_1
X_6170_ _3077_ VGND VGND VPWR VPWR _3078_ sky130_fd_sc_hd__clkbuf_1
X_5121_ tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[2\] _2125_ _0018_ VGND
+ VGND VPWR VPWR _2307_ sky130_fd_sc_hd__mux2_1
X_5052_ _0735_ _2269_ _1817_ tree_instances\[14\].u_tree.ready_for_next VGND VGND
+ VPWR VPWR _0335_ sky130_fd_sc_hd__a22o_1
X_4003_ _1471_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4743__S _0008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5954_ _2927_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5885_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[5\] VGND VGND VPWR
+ VPWR _2885_ sky130_fd_sc_hd__inv_2
X_4905_ _1641_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[5\] VGND
+ VGND VPWR VPWR _2185_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4836_ tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[3\] _1835_ _0010_ VGND
+ VGND VPWR VPWR _2127_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6506_ clknet_leaf_102_clk _0289_ net32 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_4767_ _1613_ _2030_ VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_31_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3718_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1217_ sky130_fd_sc_hd__buf_1
XTAP_TAPCELL_ROW_95_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4698_ tree_instances\[10\].u_tree.prediction_out tree_instances\[10\].u_tree.pipeline_prediction\[0\]\[0\]
+ tree_instances\[10\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6437_ clknet_leaf_23_clk _0230_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3649_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[6\] _1157_ VGND VGND
+ VPWR VPWR _1158_ sky130_fd_sc_hd__or2_1
X_6368_ clknet_leaf_19_clk _0175_ net24 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5319_ _2432_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6299_ clknet_leaf_16_clk _0108_ net29 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_59_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_39_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5670_ _2713_ tree_instances\[2\].u_tree.frame_id_out\[1\] tree_instances\[2\].u_tree.frame_id_out\[2\]
+ _2714_ VGND VGND VPWR VPWR _2715_ sky130_fd_sc_hd__o22a_1
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_32 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_0_clk_A net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4621_ _1799_ _1937_ VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__and2_1
X_4552_ _1757_ _1945_ VGND VGND VPWR VPWR _1949_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5117__A1 _2122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4483_ _1046_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[4\] VGND
+ VGND VPWR VPWR _1905_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3503_ tree_instances\[12\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__buf_1
X_3434_ _0966_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
X_6222_ _3107_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__clkbuf_1
X_3365_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _0904_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_90_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_40 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6153_ _2218_ _2171_ _3059_ _3063_ VGND VGND VPWR VPWR _3064_ sky130_fd_sc_hd__nor4_1
X_5104_ _2298_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__clkbuf_1
X_3296_ _0838_ _0840_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__nor2_1
X_6084_ _3021_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__clkbuf_1
X_5035_ _1666_ _2222_ VGND VGND VPWR VPWR _2261_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_0_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6986_ clknet_leaf_15_clk _0692_ net29 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_36_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5937_ tree_instances\[2\].u_tree.frame_id_out\[1\] tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0755_ VGND VGND VPWR VPWR _2919_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5868_ tree_instances\[1\].u_tree.frame_id_out\[0\] tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _1227_ VGND VGND VPWR VPWR _2875_ sky130_fd_sc_hd__mux2_1
X_4819_ _2117_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5799_ _2580_ _2583_ net21 VGND VGND VPWR VPWR _2837_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_8_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_2_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_19_Right_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6637__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_28_Right_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3150_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_6_Left_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_37_Right_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6840_ clknet_leaf_69_clk _0560_ net39 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6771_ clknet_leaf_5_clk _0505_ net26 VGND VGND VPWR VPWR attack_votes\[0\] sky130_fd_sc_hd__dfrtp_2
X_3983_ _1460_ _1461_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_61_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5722_ _2714_ tree_instances\[15\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2767_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_33_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6378__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5653_ attack_votes\[2\] _2700_ _2690_ VGND VGND VPWR VPWR _2701_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6307__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4604_ _1976_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5584_ _2627_ _2628_ _2629_ _2633_ VGND VGND VPWR VPWR _2634_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_46_Right_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4535_ tree_instances\[8\].u_tree.frame_id_out\[2\] tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _1000_ VGND VGND VPWR VPWR _1940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4466_ _0724_ VGND VGND VPWR VPWR _1889_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3417_ tree_instances\[11\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6205_ tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[3\] _1834_ _0036_ VGND
+ VGND VPWR VPWR _3098_ sky130_fd_sc_hd__mux2_1
X_4397_ tree_instances\[0\].u_tree.frame_id_in\[4\] VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__clkbuf_4
X_3348_ _0888_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__clkbuf_1
X_6136_ tree_instances\[17\].u_tree.pipeline_valid\[0\] tree_instances\[17\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _3049_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_55_Right_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6067_ _3009_ VGND VGND VPWR VPWR _3010_ sky130_fd_sc_hd__clkbuf_1
X_3279_ _0823_ _0825_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__or2_1
X_5018_ tree_instances\[0\].u_tree.frame_id_in\[4\] VGND VGND VPWR VPWR _2251_ sky130_fd_sc_hd__buf_4
XFILLER_0_68_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6969_ clknet_leaf_96_clk _0675_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_64_Right_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6730__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5047__B _2222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6561__SET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_73_Right_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6889__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6818__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5568__A1 _2600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_82_Right_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6471__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6400__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_10_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5740__B2 _2708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5740__A1 _2583_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4320_ _1770_ VGND VGND VPWR VPWR _1787_ sky130_fd_sc_hd__clkbuf_1
X_4251_ _1719_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_91_Right_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3202_ tree_instances\[18\].u_tree.tree_state\[0\] _0752_ _0753_ VGND VGND VPWR VPWR
+ _0063_ sky130_fd_sc_hd__a21o_1
X_4182_ _1653_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6008__S _0032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6559__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_46_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6823_ clknet_leaf_39_clk _0544_ net30 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6754_ clknet_leaf_27_clk _0008_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3966_ _1437_ VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6685_ clknet_leaf_55_clk _0434_ net35 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5705_ tree_instances\[0\].u_tree.frame_id_out\[3\] _2606_ tree_instances\[0\].u_tree.frame_id_out\[0\]
+ _2598_ VGND VGND VPWR VPWR _2750_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_57_193 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3897_ _1373_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5636_ _2659_ tree_instances\[16\].u_tree.frame_id_out\[3\] _2684_ _2685_ VGND VGND
+ VPWR VPWR _2686_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5567_ _2579_ tree_instances\[5\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2617_
+ sky130_fd_sc_hd__nor2_1
X_5498_ _2562_ VGND VGND VPWR VPWR _2563_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4518_ tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[2\] _1832_ _0042_ VGND
+ VGND VPWR VPWR _1929_ sky130_fd_sc_hd__mux2_1
X_4449_ _1876_ VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6119_ _1325_ _2972_ VGND VGND VPWR VPWR _3041_ sky130_fd_sc_hd__and2_1
XANTENNA__6982__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6911__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4836__S _0010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5521__A _2579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5789__B2 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_96_Left_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3820_ _1308_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_43_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3751_ _1242_ _1244_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6470_ clknet_leaf_29_clk _0258_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3682_ _0855_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__buf_1
X_5421_ tree_instances\[1\].u_tree.read_enable _2517_ VGND VGND VPWR VPWR _2518_ sky130_fd_sc_hd__nand2_2
XTAP_TAPCELL_ROW_76_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5352_ _2453_ VGND VGND VPWR VPWR _2454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4303_ _1765_ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5283_ tree_instances\[18\].u_tree.tree_state\[1\] tree_instances\[18\].u_tree.tree_state\[2\]
+ _1801_ VGND VGND VPWR VPWR _2413_ sky130_fd_sc_hd__or3_1
X_4234_ _0838_ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__clkbuf_1
X_4165_ _1124_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4096_ _1550_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_87_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6393__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_42_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6806_ clknet_leaf_41_clk _0528_ net36 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4998_ _1669_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[6\] _2189_
+ VGND VGND VPWR VPWR _2238_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3949_ _1412_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__clkbuf_1
X_6737_ clknet_leaf_68_clk _0485_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6668_ clknet_leaf_32_clk _0418_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6599_ clknet_leaf_60_clk _0363_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5619_ current_voting_frame\[0\] tree_instances\[12\].u_tree.frame_id_out\[0\] VGND
+ VGND VPWR VPWR _2669_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_100_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_29_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4391__S _0040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_108_Right_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5516__A _2575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5970_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[7\] tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ VGND VGND VPWR VPWR _2937_ sky130_fd_sc_hd__xor2_1
XFILLER_0_59_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4921_ _2196_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4852_ tree_instances\[12\].u_tree.frame_id_out\[3\] tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0829_ VGND VGND VPWR VPWR _2137_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_82_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_82_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3803_ _1209_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4783_ tree_instances\[12\].u_tree.tree_state\[1\] tree_instances\[12\].u_tree.current_node_data\[12\]
+ tree_instances\[12\].u_tree.node_data\[12\] _2086_ VGND VGND VPWR VPWR _2087_ sky130_fd_sc_hd__a22o_1
X_3734_ _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__clkbuf_1
X_6522_ clknet_leaf_9_clk _0305_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
X_6453_ clknet_leaf_98_clk _0246_ net26 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3665_ _1169_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload40 clknet_leaf_28_clk VGND VGND VPWR VPWR clkload40/Y sky130_fd_sc_hd__clkinv_4
Xclkload51 clknet_leaf_35_clk VGND VGND VPWR VPWR clkload51/X sky130_fd_sc_hd__clkbuf_1
XANTENNA__6021__S _0799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload62 clknet_leaf_85_clk VGND VGND VPWR VPWR clkload62/Y sky130_fd_sc_hd__inv_6
X_5404_ tree_instances\[20\].u_tree.read_enable VGND VGND VPWR VPWR _2502_ sky130_fd_sc_hd__buf_1
Xclkload84 clknet_leaf_48_clk VGND VGND VPWR VPWR clkload84/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_100_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload95 clknet_leaf_58_clk VGND VGND VPWR VPWR clkload95/Y sky130_fd_sc_hd__inv_6
X_6384_ clknet_leaf_18_clk _0191_ net24 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
Xclkload73 clknet_leaf_76_clk VGND VGND VPWR VPWR clkload73/Y sky130_fd_sc_hd__clkinvlp_4
X_3596_ _0730_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__buf_4
X_5335_ _2440_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__clkbuf_1
X_5266_ _2404_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4217_ tree_instances\[3\].u_tree.prediction_valid _0799_ VGND VGND VPWR VPWR _1688_
+ sky130_fd_sc_hd__and2b_1
X_5197_ _2326_ _2367_ VGND VGND VPWR VPWR _2369_ sky130_fd_sc_hd__and2_1
XANTENNA__6574__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4148_ _1619_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__clkbuf_1
X_4079_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1554_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6503__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_26_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_54_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5925__A1 _1829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_163 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload1 clknet_3_1__leaf_clk VGND VGND VPWR VPWR clkload1/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_34_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6102__A1 tree_instances\[0\].u_tree.frame_id_in\[4\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_69_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xload_slew35 net36 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__buf_12
XFILLER_0_84_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_111 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_37_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3450_ _0979_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3381_ _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5120_ _2306_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__clkbuf_1
X_5051_ tree_instances\[14\].u_tree.tree_state\[0\] _0734_ VGND VGND VPWR VPWR _2269_
+ sky130_fd_sc_hd__nand2_1
X_4002_ _1479_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5953_ _1421_ _2553_ VGND VGND VPWR VPWR _2927_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_51_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4904_ _0958_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[1\] VGND
+ VGND VPWR VPWR _2184_ sky130_fd_sc_hd__and2b_1
XTAP_TAPCELL_ROW_23_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5884_ _1394_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[6\] _2883_
+ VGND VGND VPWR VPWR _2884_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4835_ _2126_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4766_ _2078_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__clkbuf_1
X_3717_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1216_ sky130_fd_sc_hd__buf_1
X_6505_ clknet_leaf_101_clk _0288_ net32 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_31_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_95_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4697_ _2035_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__clkbuf_1
X_6436_ clknet_leaf_18_clk _0229_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3648_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1157_ sky130_fd_sc_hd__buf_1
XFILLER_0_3_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3579_ _1096_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__clkbuf_1
X_6367_ clknet_leaf_19_clk _0174_ net24 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6755__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5318_ tree_instances\[19\].u_tree.frame_id_out\[4\] tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[19\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2432_ sky130_fd_sc_hd__mux2_1
X_6298_ _0903_ _3148_ _0036_ tree_instances\[5\].u_tree.pipeline_valid\[0\] VGND VGND
+ VPWR VPWR _0704_ sky130_fd_sc_hd__o2bb2a_1
X_5249_ _2395_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6425__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkload4_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4620_ _1984_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4551_ _1948_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3502_ tree_instances\[9\].u_tree.tree_state\[0\] _1024_ _1025_ VGND VGND VPWR VPWR
+ _0085_ sky130_fd_sc_hd__a21o_1
X_4482_ _1765_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[3\] VGND
+ VGND VPWR VPWR _1904_ sky130_fd_sc_hd__or2_1
X_3433_ _0965_ tree_instances\[13\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0966_
+ sky130_fd_sc_hd__and2b_1
X_6221_ tree_instances\[5\].u_tree.frame_id_out\[4\] tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[5\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _3107_ sky130_fd_sc_hd__mux2_1
X_6152_ _2175_ _3062_ _2182_ _2172_ VGND VGND VPWR VPWR _3063_ sky130_fd_sc_hd__or4b_1
X_5103_ _1455_ _2296_ VGND VGND VPWR VPWR _2298_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3364_ tree_instances\[5\].u_tree.tree_state\[0\] _0902_ _0903_ VGND VGND VPWR VPWR
+ _0077_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_90_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__buf_1
X_6083_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[4\] _1344_ _3020_
+ VGND VGND VPWR VPWR _3021_ sky130_fd_sc_hd__mux2_1
X_5034_ _2260_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_0_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6985_ clknet_leaf_38_clk _0691_ net30 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5053__A1 _2122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_64_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5936_ _2918_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__clkbuf_1
X_5867_ _2873_ _2874_ _2534_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4818_ _1278_ _2071_ VGND VGND VPWR VPWR _2117_ sky130_fd_sc_hd__and2_1
X_5798_ _2713_ net21 VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4749_ tree_instances\[10\].u_tree.current_node_data\[12\] tree_instances\[10\].u_tree.node_data\[12\]
+ _1172_ VGND VGND VPWR VPWR _2069_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6936__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6419_ clknet_leaf_57_clk _0064_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6677__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6606__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3982_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1461_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6770_ clknet_leaf_11_clk _0504_ net29 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.frame_id_in\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_43_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5721_ _2708_ tree_instances\[15\].u_tree.frame_id_out\[4\] _2765_ VGND VGND VPWR
+ VPWR _2766_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_61_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5652_ _2572_ _2699_ VGND VGND VPWR VPWR _2700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4603_ tree_instances\[9\].u_tree.frame_id_out\[1\] tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _1025_ VGND VGND VPWR VPWR _1976_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5583_ _2579_ _2630_ tree_instances\[3\].u_tree.frame_id_out\[4\] _2631_ _2632_ VGND
+ VGND VPWR VPWR _2633_ sky130_fd_sc_hd__o221a_1
XFILLER_0_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_107_Left_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4534_ _1939_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6347__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4465_ _1887_ VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4396_ _1836_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
X_3416_ _0934_ _0943_ _0947_ _0950_ tree_instances\[5\].u_tree.tree_state\[1\] VGND
+ VGND VPWR VPWR _0078_ sky130_fd_sc_hd__a41o_1
X_6204_ _3097_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__clkbuf_1
X_3347_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _0888_ sky130_fd_sc_hd__inv_2
X_6135_ _0849_ _1955_ _1807_ tree_instances\[4\].u_tree.ready_for_next VGND VGND VPWR
+ VPWR _0641_ sky130_fd_sc_hd__a22o_1
X_6066_ _3008_ VGND VGND VPWR VPWR _3009_ sky130_fd_sc_hd__clkbuf_1
X_5017_ _2250_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__clkbuf_1
X_3278_ _0824_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_101_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6968_ clknet_leaf_81_clk _0674_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_6899_ clknet_leaf_33_clk _0001_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.gen_tree_16.u_tree_rom.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6657__SET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5919_ _2152_ _2900_ VGND VGND VPWR VPWR _2910_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6770__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_67_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6858__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_10_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6440__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4250_ _1710_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3201_ tree_instances\[18\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__buf_2
X_4181_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1653_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5008__A1 _2122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6822_ clknet_leaf_39_clk _0543_ net30 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_18_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6753_ clknet_leaf_27_clk _0007_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3965_ _1440_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3896_ _1367_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__clkbuf_1
X_6684_ clknet_leaf_56_clk _0433_ net35 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5704_ tree_instances\[0\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2749_ sky130_fd_sc_hd__inv_2
XANTENNA__6599__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5635_ tree_instances\[16\].u_tree.frame_id_out\[1\] _2579_ VGND VGND VPWR VPWR _2685_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__6528__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5566_ _2578_ tree_instances\[5\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2616_
+ sky130_fd_sc_hd__and2_1
X_5497_ _0725_ VGND VGND VPWR VPWR _2562_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4517_ _1928_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4448_ _1875_ VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5615__A_N _2585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4379_ _1824_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__inv_2
X_6118_ _3040_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__clkbuf_1
X_6049_ _2450_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[1\] _2990_
+ _2991_ tree_instances\[5\].u_tree.u_tree_weight_rom.cache_valid VGND VGND VPWR VPWR
+ _2992_ sky130_fd_sc_hd__o221a_1
XFILLER_0_64_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6951__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5802__A _2586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6692__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3750_ _1243_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3681_ _1185_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5420_ _1496_ _2504_ _2510_ _2511_ _2516_ VGND VGND VPWR VPWR _2517_ sky130_fd_sc_hd__a2111o_1
XTAP_TAPCELL_ROW_76_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_9 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5351_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _2453_ sky130_fd_sc_hd__inv_2
X_5282_ _2412_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__clkbuf_1
X_4302_ _1042_ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4233_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1702_ sky130_fd_sc_hd__inv_2
X_4164_ _1628_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__clkbuf_1
X_4095_ _1565_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_87_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6805_ clknet_leaf_41_clk _0527_ net36 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_91 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6736_ clknet_leaf_67_clk _0484_ net36 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4997_ _2237_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_621 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3948_ _1427_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3879_ _1361_ _1362_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__nor2_1
X_6667_ clknet_leaf_30_clk _0417_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_21_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6598_ clknet_leaf_60_clk _0362_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5618_ tree_instances\[12\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2668_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5549_ _2582_ VGND VGND VPWR VPWR _2599_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_29_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4920_ _1724_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[3\] _2192_
+ VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6802__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4851_ _2136_ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_82_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3802_ _1212_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5395__B1 _0004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4782_ tree_instances\[12\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _2086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3733_ _1229_ _0898_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6521_ clknet_leaf_8_clk _0304_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.prediction_out
+ sky130_fd_sc_hd__dfrtp_1
X_6452_ clknet_leaf_98_clk _0245_ net26 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3664_ _1171_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__buf_1
XFILLER_0_43_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload41 clknet_leaf_29_clk VGND VGND VPWR VPWR clkload41/X sky130_fd_sc_hd__clkbuf_1
Xclkload52 clknet_leaf_36_clk VGND VGND VPWR VPWR clkload52/Y sky130_fd_sc_hd__clkinv_2
Xclkload30 clknet_leaf_17_clk VGND VGND VPWR VPWR clkload30/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5403_ _2501_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__clkbuf_1
Xclkload85 clknet_leaf_49_clk VGND VGND VPWR VPWR clkload85/Y sky130_fd_sc_hd__clkinv_4
Xclkload96 clknet_leaf_59_clk VGND VGND VPWR VPWR clkload96/Y sky130_fd_sc_hd__bufinv_16
Xclkload74 clknet_leaf_77_clk VGND VGND VPWR VPWR clkload74/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6383_ clknet_leaf_84_clk _0190_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[7\] sky130_fd_sc_hd__dfrtp_1
X_3595_ _1108_ _1111_ tree_instances\[8\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR
+ _0041_ sky130_fd_sc_hd__o21a_1
Xclkload63 clknet_leaf_86_clk VGND VGND VPWR VPWR clkload63/Y sky130_fd_sc_hd__bufinv_16
X_5334_ _1561_ _2413_ VGND VGND VPWR VPWR _2440_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5265_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[4\] _1380_ _2399_
+ VGND VGND VPWR VPWR _2404_ sky130_fd_sc_hd__mux2_1
X_5196_ _2368_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__clkbuf_1
X_4216_ _1687_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4147_ tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4078_ _1551_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5622__B2 tree_instances\[12\].u_tree.prediction_out VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__6543__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_440 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6719_ clknet_leaf_47_clk _0467_ net34 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload2 clknet_3_3__leaf_clk VGND VGND VPWR VPWR clkload2/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5689__A1 _2622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5689__B2 _2631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xload_slew36 net39 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__buf_12
XFILLER_0_96_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_3_4__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3380_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__7001__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_41_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5050_ _2268_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__clkbuf_1
X_4001_ _1478_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_56_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5952_ _2926_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5604__B2 _2619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5604__A1 _2576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4903_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[1\] _0958_ VGND
+ VGND VPWR VPWR _2183_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5883_ _1404_ _2881_ _2882_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[7\]
+ VGND VGND VPWR VPWR _2883_ sky130_fd_sc_hd__a22o_1
X_4834_ tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[2\] _2125_ _0010_ VGND
+ VGND VPWR VPWR _2126_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4765_ _1607_ _2030_ VGND VGND VPWR VPWR _2078_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3716_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[7\] _0914_ VGND VGND
+ VPWR VPWR _1215_ sky130_fd_sc_hd__or2_1
XANTENNA__4591__A1 _1830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6504_ clknet_leaf_100_clk _0287_ net32 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_95_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4696_ tree_instances\[10\].u_tree.frame_id_out\[4\] tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[10\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_31_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3647_ _1140_ _1148_ _1153_ _1156_ tree_instances\[11\].u_tree.tree_state\[1\] VGND
+ VGND VPWR VPWR _0050_ sky130_fd_sc_hd__a41o_1
X_6435_ clknet_leaf_18_clk _0228_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6366_ clknet_leaf_15_clk _0173_ net29 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3578_ _1095_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5317_ _2431_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6096__A1 _1829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6297_ tree_instances\[5\].u_tree.pipeline_valid\[0\] tree_instances\[5\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _3148_ sky130_fd_sc_hd__nand2_1
X_5248_ _1388_ _2314_ VGND VGND VPWR VPWR _2395_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_59_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5179_ _1217_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND
+ VGND VPWR VPWR _2353_ sky130_fd_sc_hd__nor2_1
XANTENNA__6795__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6724__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_3_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_39_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6465__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4550_ _1760_ _1945_ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3501_ tree_instances\[9\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__buf_2
X_4481_ _1770_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[3\] VGND
+ VGND VPWR VPWR _1903_ sky130_fd_sc_hd__nand2_1
XANTENNA__5522__A0 _2580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3432_ _0955_ _0961_ _0964_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__and3b_1
X_6220_ _3106_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6151_ _3060_ _3061_ _2178_ _2185_ VGND VGND VPWR VPWR _3062_ sky130_fd_sc_hd__or4_1
X_3363_ tree_instances\[5\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__buf_2
X_5102_ _2297_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_29_Left_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_90_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0839_ sky130_fd_sc_hd__buf_1
X_6082_ _2988_ VGND VGND VPWR VPWR _3020_ sky130_fd_sc_hd__clkbuf_2
X_5033_ tree_instances\[14\].u_tree.frame_id_out\[4\] tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[14\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2260_ sky130_fd_sc_hd__mux2_1
XANTENNA__6027__S _0799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6984_ clknet_leaf_16_clk _0690_ net29 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_64_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5935_ tree_instances\[2\].u_tree.frame_id_out\[0\] tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0755_ VGND VGND VPWR VPWR _2918_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_36_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5866_ tree_instances\[1\].u_tree.tree_state\[1\] _2856_ VGND VGND VPWR VPWR _2874_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_38_Left_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4817_ _2116_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_131 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5797_ net21 _2836_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4748_ _2068_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4679_ _2024_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6418_ clknet_leaf_56_clk _0022_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_1_Right_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_8_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6349_ clknet_leaf_21_clk _0156_ net24 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6617__SET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5630__A _2610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6646__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5807__A1 _1826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3981_ _1459_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5720_ _2708_ tree_instances\[15\].u_tree.frame_id_out\[4\] tree_instances\[15\].u_tree.frame_id_out\[3\]
+ _2709_ VGND VGND VPWR VPWR _2765_ sky130_fd_sc_hd__a2bb2o_1
XTAP_TAPCELL_ROW_61_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_33_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_42_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5651_ attack_votes\[0\] attack_votes\[1\] attack_votes\[2\] VGND VGND VPWR VPWR
+ _2699_ sky130_fd_sc_hd__and3_1
X_4602_ _1975_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
X_5582_ _2582_ tree_instances\[3\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2632_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_13_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4533_ tree_instances\[8\].u_tree.frame_id_out\[1\] tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _1000_ VGND VGND VPWR VPWR _1939_ sky130_fd_sc_hd__mux2_1
XANTENNA__5715__A _2588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4464_ _1886_ VGND VGND VPWR VPWR _1887_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6203_ tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[2\] _2595_ _0036_ VGND
+ VGND VPWR VPWR _3097_ sky130_fd_sc_hd__mux2_1
XFILLER_0_68_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4395_ tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[3\] _1835_ _0040_ VGND
+ VGND VPWR VPWR _1836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3415_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[6\] _0949_ VGND VGND
+ VPWR VPWR _0950_ sky130_fd_sc_hd__nor2_1
X_3346_ _0886_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__clkbuf_1
X_6134_ _3048_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6316__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6065_ net42 VGND VGND VPWR VPWR _3008_ sky130_fd_sc_hd__clkbuf_1
X_5016_ tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[3\] _2249_ _0014_ VGND
+ VGND VPWR VPWR _2250_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3277_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _0824_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6967_ clknet_leaf_96_clk _0673_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_101_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5918_ _2909_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_33_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6898_ clknet_leaf_83_clk _0612_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.node_data\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5849_ _2864_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_110 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_24_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_10_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6827__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3200_ _0733_ tree_instances\[18\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _0752_ sky130_fd_sc_hd__or2_1
X_4180_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1652_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6480__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6821_ clknet_leaf_39_clk _0542_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6205__A1 _1834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_46_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6752_ clknet_leaf_24_clk _0049_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
Xclkbuf_leaf_15_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_4
X_3964_ _1443_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3895_ _1371_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__clkbuf_1
X_6683_ clknet_leaf_44_clk _0432_ net34 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5703_ _2746_ _2583_ tree_instances\[0\].u_tree.frame_id_out\[3\] _2659_ _2747_ VGND
+ VGND VPWR VPWR _2748_ sky130_fd_sc_hd__o221a_1
X_5634_ _2578_ tree_instances\[16\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2684_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_232 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5565_ _2588_ tree_instances\[5\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2615_
+ sky130_fd_sc_hd__xnor2_1
X_5496_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[8\] VGND VGND VPWR
+ VPWR _2561_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6568__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4516_ tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[1\] _1830_ _0042_ VGND
+ VGND VPWR VPWR _1928_ sky130_fd_sc_hd__mux2_1
X_4447_ _1874_ VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6117_ tree_instances\[4\].u_tree.frame_id_out\[4\] tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[4\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _3040_ sky130_fd_sc_hd__mux2_1
X_4378_ _1823_ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__buf_2
X_3329_ _0870_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__clkbuf_1
X_6048_ _0937_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[3\] VGND
+ VGND VPWR VPWR _2991_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6991__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6920__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_73_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_43_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3680_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[5\] _0852_ VGND VGND
+ VPWR VPWR _1185_ sky130_fd_sc_hd__or2_1
XFILLER_0_23_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5350_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _2452_ sky130_fd_sc_hd__clkbuf_1
X_5281_ tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[4\] _2251_ _0022_ VGND
+ VGND VPWR VPWR _2412_ sky130_fd_sc_hd__mux2_1
XFILLER_0_64_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4301_ _1767_ VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4232_ _1700_ VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_4_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_4
X_4163_ _1629_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4094_ _1256_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_87_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_63 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6804_ clknet_leaf_42_clk _0526_ net36 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4996_ _1676_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[5\] _2189_
+ VGND VGND VPWR VPWR _2237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_238 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3947_ _0758_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__clkbuf_1
X_6735_ clknet_leaf_68_clk _0483_ net36 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6666_ clknet_leaf_29_clk _0416_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_3878_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[7\] tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[6\]
+ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6749__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6597_ clknet_leaf_59_clk _0361_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5617_ _2603_ tree_instances\[12\].u_tree.frame_id_out\[1\] _2665_ _2666_ VGND VGND
+ VPWR VPWR _2667_ sky130_fd_sc_hd__a211oi_1
X_5548_ _2575_ VGND VGND VPWR VPWR _2598_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6331__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5479_ _2552_ VGND VGND VPWR VPWR _2553_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_29_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_107_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6419__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_0_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4850_ tree_instances\[12\].u_tree.frame_id_out\[2\] tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0829_ VGND VGND VPWR VPWR _2136_ sky130_fd_sc_hd__mux2_1
X_3801_ _1289_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4781_ _2085_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__clkbuf_1
X_6520_ clknet_leaf_8_clk _0303_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3732_ _0897_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6842__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5707__B _2579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6451_ clknet_leaf_97_clk _0244_ net32 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4611__B _1937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3663_ tree_instances\[10\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload20 clknet_leaf_10_clk VGND VGND VPWR VPWR clkload20/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload42 clknet_leaf_30_clk VGND VGND VPWR VPWR clkload42/Y sky130_fd_sc_hd__clkinv_1
Xclkload53 clknet_leaf_37_clk VGND VGND VPWR VPWR clkload53/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload31 clknet_leaf_18_clk VGND VGND VPWR VPWR clkload31/Y sky130_fd_sc_hd__clkinvlp_4
X_6382_ clknet_leaf_79_clk _0189_ net39 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_5402_ tree_instances\[20\].u_tree.pipeline_prediction\[0\]\[0\] _2498_ _2500_ VGND
+ VGND VPWR VPWR _2501_ sky130_fd_sc_hd__mux2_1
Xclkload86 clknet_leaf_50_clk VGND VGND VPWR VPWR clkload86/Y sky130_fd_sc_hd__bufinv_16
X_5333_ _2439_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__clkbuf_1
Xclkload75 clknet_leaf_78_clk VGND VGND VPWR VPWR clkload75/Y sky130_fd_sc_hd__clkinvlp_4
X_3594_ _1110_ _1045_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload64 clknet_leaf_87_clk VGND VGND VPWR VPWR clkload64/Y sky130_fd_sc_hd__bufinv_16
XFILLER_0_100_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload97 clknet_leaf_60_clk VGND VGND VPWR VPWR clkload97/Y sky130_fd_sc_hd__bufinv_16
XPHY_EDGE_ROW_10_Left_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5264_ _2403_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__clkbuf_1
X_5195_ _2325_ _2367_ VGND VGND VPWR VPWR _2368_ sky130_fd_sc_hd__and2_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4215_ tree_instances\[2\].u_tree.prediction_valid _0755_ VGND VGND VPWR VPWR _1687_
+ sky130_fd_sc_hd__and2b_1
X_7003_ clknet_leaf_87_clk _0704_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4146_ _1618_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4077_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_54_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4979_ tree_instances\[13\].u_tree.prediction_out tree_instances\[13\].u_tree.pipeline_prediction\[0\]\[0\]
+ tree_instances\[13\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_452 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6583__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6718_ clknet_leaf_48_clk _0466_ net34 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload3 clknet_3_4__leaf_clk VGND VGND VPWR VPWR clkload3/X sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6649_ clknet_leaf_31_clk _0408_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6512__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5633__A _2622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_70_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew37 net38 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_12
XFILLER_0_69_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4000_ _1477_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5951_ _1432_ _2553_ VGND VGND VPWR VPWR _2926_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4902_ _1656_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND
+ VGND VPWR VPWR _2182_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_51_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5882_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[7\] VGND VGND VPWR
+ VPWR _2882_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4833_ tree_instances\[0\].u_tree.frame_id_in\[2\] VGND VGND VPWR VPWR _2125_ sky130_fd_sc_hd__buf_4
X_4764_ _2077_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3715_ _1207_ _1208_ _1214_ _1001_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__o31a_1
X_6503_ clknet_leaf_101_clk _0286_ net32 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6434_ clknet_leaf_95_clk _0227_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.cached_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4695_ _2034_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__clkbuf_1
X_3646_ _1154_ _1155_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_95_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3577_ _1093_ _1094_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6365_ clknet_leaf_11_clk _0172_ net29 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6296_ _0932_ _3081_ _1811_ tree_instances\[6\].u_tree.ready_for_next VGND VGND VPWR
+ VPWR _0703_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5316_ tree_instances\[19\].u_tree.frame_id_out\[3\] tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _1252_ VGND VGND VPWR VPWR _2431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5247_ _2394_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_59_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5178_ _1375_ _2348_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ _1355_ _2351_ VGND VGND VPWR VPWR _2352_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_3_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4129_ _1603_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_104_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6764__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_load_slew35_A net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5598__A1 _2598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5598__B2 _2606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6928__SET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5770__B2 _2603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5770__A1 _2598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3500_ _0733_ tree_instances\[9\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _1024_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4480_ _1901_ VGND VGND VPWR VPWR _1902_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3431_ _0963_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6150_ _1658_ _2170_ _2173_ VGND VGND VPWR VPWR _3061_ sky130_fd_sc_hd__o21ai_1
X_3362_ _0732_ tree_instances\[5\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _0902_ sky130_fd_sc_hd__or2_1
X_5101_ _1442_ _2296_ VGND VGND VPWR VPWR _2297_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_182 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_90_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3293_ _0837_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__buf_1
X_6081_ _3019_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__clkbuf_1
X_5032_ _2259_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_0_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6983_ clknet_leaf_38_clk _0689_ net30 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_0_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_64_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5934_ _2917_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__clkbuf_1
X_5865_ _2872_ VGND VGND VPWR VPWR _2873_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4816_ _1274_ _2071_ VGND VGND VPWR VPWR _2116_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4352__A _1803_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5796_ _2627_ _0000_ VGND VGND VPWR VPWR _2836_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4747_ tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[4\] _1837_ _0008_ VGND
+ VGND VPWR VPWR _2068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5761__B2 _2708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5761__A1 _2603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_444 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4678_ tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[3\] _1835_ _0006_ VGND
+ VGND VPWR VPWR _2024_ sky130_fd_sc_hd__mux2_1
X_6417_ clknet_leaf_56_clk _0021_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3629_ _1139_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6348_ clknet_leaf_20_clk _0155_ net26 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_8_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6279_ _3139_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6945__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_40_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5752__A1 _2583_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_55_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6686__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6615__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3980_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1459_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_61_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_0_clk net40 VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_5650_ _1018_ _2696_ _2697_ _2698_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__a31o_1
X_4601_ tree_instances\[9\].u_tree.frame_id_out\[0\] tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _1025_ VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__mux2_1
XANTENNA__5743__A1 _2586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5581_ current_voting_frame\[4\] VGND VGND VPWR VPWR _2631_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_13_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4532_ _1938_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
X_4463_ _0716_ VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3414_ _0948_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__clkbuf_1
X_6202_ _3096_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_15_Right_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4394_ _1834_ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__clkbuf_4
X_3345_ _0884_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__or2_1
X_6133_ _1346_ _2971_ VGND VGND VPWR VPWR _3048_ sky130_fd_sc_hd__and2_1
X_6064_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[7\] _2489_ _3005_ _3006_
+ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[8\] VGND VGND VPWR VPWR _3007_
+ sky130_fd_sc_hd__a2111oi_1
X_3276_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _0823_ sky130_fd_sc_hd__clkbuf_1
X_5015_ tree_instances\[0\].u_tree.frame_id_in\[3\] VGND VGND VPWR VPWR _2249_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6966_ clknet_leaf_46_clk _0002_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.gen_tree_1.u_tree_rom.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XPHY_EDGE_ROW_24_Right_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_101_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5917_ _2159_ _2900_ VGND VGND VPWR VPWR _2909_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6897_ clknet_leaf_70_clk _0611_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.node_data\[107\]
+ sky130_fd_sc_hd__dfxtp_1
X_5848_ _1525_ _2427_ VGND VGND VPWR VPWR _2864_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5734__A1 _2709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5779_ complete_votes\[1\] VGND VGND VPWR VPWR _2823_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_2_Left_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_33_Right_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_42_Right_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5725__B2 _2709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5725__A1 _2713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_57_Left_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_51_Right_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_78_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6867__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_66_Left_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_60_Right_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6820_ clknet_leaf_55_clk _0541_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_18_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3963_ _1052_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6751_ clknet_leaf_92_clk _0048_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3894_ _1370_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__clkbuf_1
X_6682_ clknet_leaf_51_clk _0431_ net35 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5702_ tree_instances\[0\].u_tree.frame_id_out\[4\] _2588_ VGND VGND VPWR VPWR _2747_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_75_Left_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5633_ _2622_ tree_instances\[16\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2683_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__5716__A1 _2606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5564_ tree_instances\[20\].u_tree.prediction_out _2613_ VGND VGND VPWR VPWR _2614_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_79_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4515_ _1927_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_103_Right_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5495_ _1023_ _2560_ _0018_ tree_instances\[16\].u_tree.pipeline_valid\[0\] VGND
+ VGND VPWR VPWR _0488_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_13_244 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4446_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1874_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4377_ _1822_ _1113_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__or2_1
X_3328_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _0870_ sky130_fd_sc_hd__clkbuf_1
X_6116_ _3039_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_84_Left_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6047_ _2452_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[3\] VGND
+ VGND VPWR VPWR _2990_ sky130_fd_sc_hd__and2_1
X_3259_ _0804_ _0805_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6949_ clknet_leaf_87_clk _0661_ net30 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_73_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6960__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6199__A1 _1826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_max_cap39_A tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_43_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5546__A _1837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_328 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5280_ _2411_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__clkbuf_1
X_4300_ _1041_ _1766_ VGND VGND VPWR VPWR _1767_ sky130_fd_sc_hd__or2_1
XANTENNA__6454__SET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4231_ _1692_ _1694_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__nor2_1
XFILLER_0_49_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4162_ _1632_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6630__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4093_ _1553_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6803_ clknet_leaf_40_clk _0525_ net36 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4995_ _2236_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6734_ clknet_leaf_67_clk _0482_ net36 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3946_ _1416_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3877_ _1360_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__clkbuf_1
X_6665_ clknet_leaf_29_clk _0415_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_61_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_205 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_98_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6596_ clknet_leaf_59_clk _0360_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4360__A _1112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5616_ tree_instances\[12\].u_tree.frame_id_out\[3\] _2585_ VGND VGND VPWR VPWR _2666_
+ sky130_fd_sc_hd__and2b_1
XANTENNA__6742__SET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6789__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5547_ attack_votes\[0\] _1020_ VGND VGND VPWR VPWR _2597_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5478_ _0756_ tree_instances\[20\].u_tree.tree_state\[1\] _2550_ VGND VGND VPWR VPWR
+ _2552_ sky130_fd_sc_hd__or3_1
X_4429_ _0981_ VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6718__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_92_Left_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4676__A1 _1832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6371__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6300__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_107_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_40_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6459__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_56_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3800_ _1014_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4780_ _1429_ _1430_ VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__and2_1
X_3731_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6450_ clknet_leaf_97_clk _0243_ net32 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3662_ _1170_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__inv_2
Xclkload10 clknet_leaf_4_clk VGND VGND VPWR VPWR clkload10/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_70_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload32 clknet_leaf_19_clk VGND VGND VPWR VPWR clkload32/X sky130_fd_sc_hd__clkbuf_1
Xclkload43 clknet_leaf_13_clk VGND VGND VPWR VPWR clkload43/Y sky130_fd_sc_hd__clkinv_4
Xclkload21 clknet_leaf_11_clk VGND VGND VPWR VPWR clkload21/Y sky130_fd_sc_hd__clkinv_2
X_6381_ clknet_leaf_77_clk _0188_ net39 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3593_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__clkbuf_1
X_5401_ _0027_ _1198_ _2499_ VGND VGND VPWR VPWR _2500_ sky130_fd_sc_hd__and3b_1
X_5332_ _1564_ _2414_ VGND VGND VPWR VPWR _2439_ sky130_fd_sc_hd__and2_1
Xclkload54 clknet_leaf_38_clk VGND VGND VPWR VPWR clkload54/Y sky130_fd_sc_hd__clkinv_2
Xclkload87 clknet_leaf_64_clk VGND VGND VPWR VPWR clkload87/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload76 clknet_leaf_79_clk VGND VGND VPWR VPWR clkload76/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__6882__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload65 clknet_leaf_88_clk VGND VGND VPWR VPWR clkload65/Y sky130_fd_sc_hd__inv_6
XANTENNA__6811__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload98 clknet_leaf_61_clk VGND VGND VPWR VPWR clkload98/X sky130_fd_sc_hd__clkbuf_1
X_5263_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[3\] _1384_ _2399_
+ VGND VGND VPWR VPWR _2403_ sky130_fd_sc_hd__mux2_1
X_7002_ clknet_leaf_52_clk _0066_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5194_ _2366_ VGND VGND VPWR VPWR _2367_ sky130_fd_sc_hd__clkbuf_2
X_4214_ _1678_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__buf_1
XFILLER_0_76_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4145_ tree_instances\[1\].u_tree.prediction_valid _1227_ VGND VGND VPWR VPWR _1618_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4076_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_122 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4978_ _2227_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__clkbuf_1
X_6717_ clknet_leaf_35_clk _0465_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.cached_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3929_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1409_ sky130_fd_sc_hd__inv_2
Xclkload4 clknet_3_5__leaf_clk VGND VGND VPWR VPWR clkload4/Y sky130_fd_sc_hd__clkinvlp_2
XFILLER_0_34_615 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6648_ clknet_leaf_31_clk _0407_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_136 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6579_ clknet_leaf_52_clk _0348_ net35 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6552__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xload_slew38 net39 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_12
XFILLER_0_69_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5950_ _2925_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4901_ _1662_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[6\] _2178_
+ _2180_ VGND VGND VPWR VPWR _2181_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5881_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[1\] VGND VGND VPWR
+ VPWR _2881_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4832_ _2124_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4763_ _1591_ _2030_ VGND VGND VPWR VPWR _2077_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3714_ _1211_ _1213_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__nand2_1
X_6502_ clknet_leaf_102_clk _0285_ net32 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4694_ tree_instances\[10\].u_tree.frame_id_out\[3\] tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _1136_ VGND VGND VPWR VPWR _2034_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6433_ clknet_leaf_98_clk _0226_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3645_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3576_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6364_ clknet_leaf_84_clk _0171_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.cached_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_5315_ _2430_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6295_ _3147_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__clkbuf_1
X_5246_ _1383_ _2314_ VGND VGND VPWR VPWR _2394_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_89_Right_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_59_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5177_ _1367_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[1\] VGND
+ VGND VPWR VPWR _2351_ sky130_fd_sc_hd__xor2_1
X_4128_ _1157_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__clkbuf_1
X_4059_ _1086_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_3_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_39_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_98_Right_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6733__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5745__A_N _2580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_load_slew28_A net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_37 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6474__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6403__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_426 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3430_ _0962_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__clkbuf_1
X_3361_ _0895_ _0900_ _0901_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__o21a_1
XFILLER_0_0_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5100_ tree_instances\[15\].u_tree.tree_state\[2\] tree_instances\[15\].u_tree.tree_state\[1\]
+ _2275_ VGND VGND VPWR VPWR _2296_ sky130_fd_sc_hd__or3_2
XFILLER_0_0_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6080_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[3\] _1347_ _2989_
+ VGND VGND VPWR VPWR _3019_ sky130_fd_sc_hd__mux2_1
X_5031_ tree_instances\[14\].u_tree.frame_id_out\[3\] tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0735_ VGND VGND VPWR VPWR _2259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3292_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _0837_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4617__B _1937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_0_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6982_ clknet_leaf_83_clk _0688_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.current_node_data\[107\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_64_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5933_ tree_instances\[20\].u_tree.current_node_data\[12\] tree_instances\[20\].u_tree.node_data\[12\]
+ _0757_ VGND VGND VPWR VPWR _2917_ sky130_fd_sc_hd__mux2_1
X_5864_ tree_instances\[1\].u_tree.read_enable VGND VGND VPWR VPWR _2872_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4815_ _2115_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5795_ _2835_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4746_ _2067_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4677_ _2023_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6416_ clknet_leaf_62_clk _0063_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_3628_ _1137_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__or2_1
X_6347_ clknet_leaf_20_clk _0154_ net26 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_8_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3559_ _1078_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_8_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5277__A1 _2125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6278_ _2456_ _3102_ VGND VGND VPWR VPWR _3139_ sky130_fd_sc_hd__and2_1
XANTENNA__6997__SET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5229_ _2385_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6985__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6914__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkload2_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6655__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_33_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5549__A _2582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4600_ _1974_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5580_ tree_instances\[3\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2630_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_13_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4531_ tree_instances\[8\].u_tree.frame_id_out\[0\] tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _1000_ VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__mux2_1
XANTENNA__4951__A0 _1827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4462_ _0713_ VGND VGND VPWR VPWR _1885_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3413_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[4\] tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[5\]
+ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__or2_1
X_6201_ tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[1\] _1829_ _0036_ VGND
+ VGND VPWR VPWR _3096_ sky130_fd_sc_hd__mux2_1
X_4393_ tree_instances\[0\].u_tree.frame_id_in\[3\] VGND VGND VPWR VPWR _1834_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3344_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _0885_ sky130_fd_sc_hd__clkbuf_1
X_6132_ _3047_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__clkbuf_1
X_6063_ _1248_ _2483_ _2485_ _2492_ VGND VGND VPWR VPWR _3006_ sky130_fd_sc_hd__and4_1
X_3275_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[1\] _0821_ VGND VGND
+ VPWR VPWR _0822_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5014_ _2248_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6965_ clknet_leaf_50_clk _0056_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_101_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5916_ _2908_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6396__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6896_ clknet_leaf_35_clk _0610_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_5847_ _2863_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6325__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5778_ _2447_ _2707_ _2821_ _2822_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__o31a_1
X_4729_ _1608_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[4\] _2010_
+ VGND VGND VPWR VPWR _2059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_191 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5670__B2 _2714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5670__A1 _2713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_103_Left_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_98_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_67_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_101_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5646__B1_N _2636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6836__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6750_ clknet_leaf_92_clk _0006_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_46_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5701_ tree_instances\[0\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2746_ sky130_fd_sc_hd__inv_2
X_3962_ _1441_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3893_ _0913_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__clkbuf_1
X_6681_ clknet_leaf_61_clk _0430_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5632_ _2606_ tree_instances\[16\].u_tree.frame_id_out\[3\] _2680_ _2681_ tree_instances\[16\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2682_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5563_ _2601_ _2604_ _2607_ _2612_ VGND VGND VPWR VPWR _2613_ sky130_fd_sc_hd__and4_1
XFILLER_0_79_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4514_ tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[0\] _1827_ _0042_ VGND
+ VGND VPWR VPWR _1927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5494_ tree_instances\[16\].u_tree.pipeline_valid\[0\] tree_instances\[16\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _2560_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4445_ _1873_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4376_ tree_instances\[13\].u_tree.tree_state\[0\] VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__inv_2
X_3327_ _0867_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__or2_1
X_6115_ tree_instances\[4\].u_tree.frame_id_out\[3\] tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0849_ VGND VGND VPWR VPWR _3039_ sky130_fd_sc_hd__mux2_1
XANTENNA__4358__A _1803_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3258_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[5\] tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[4\]
+ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__nand2_1
X_6046_ _2988_ VGND VGND VPWR VPWR _2989_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__6577__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3189_ _0739_ _0741_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_54_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_643 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6506__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6948_ clknet_leaf_88_clk _0660_ net30 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6879_ clknet_leaf_12_clk _0598_ net29 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_69_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4391__A1 _1832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_226 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_543 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4230_ _0834_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__clkbuf_1
X_4161_ _1624_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4092_ _1552_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6670__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6802_ clknet_leaf_45_clk _0524_ net34 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4344__C net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4994_ _1647_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[4\] _2189_
+ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3945_ _1417_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__clkbuf_1
X_6733_ clknet_leaf_68_clk _0481_ net36 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6664_ clknet_leaf_33_clk _0414_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3876_ _0925_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__clkbuf_1
X_5615_ _2585_ tree_instances\[12\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2665_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6595_ clknet_leaf_60_clk _0359_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5546_ _1837_ _2596_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5477_ tree_instances\[20\].u_tree.tree_state\[1\] _2499_ VGND VGND VPWR VPWR _2551_
+ sky130_fd_sc_hd__or2b_1
X_4428_ _1859_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6758__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4359_ _1813_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__inv_2
X_6029_ tree_instances\[3\].u_tree.frame_id_out\[4\] tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[3\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2977_ sky130_fd_sc_hd__mux2_1
XANTENNA__5625__B2 _2603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5625__A1 _2598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6340__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_86_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_28_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3730_ tree_instances\[1\].u_tree.tree_state\[0\] _1226_ _1227_ VGND VGND VPWR VPWR
+ _0067_ sky130_fd_sc_hd__a21o_1
XFILLER_0_67_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3661_ tree_instances\[10\].u_tree.tree_state\[2\] _1169_ VGND VGND VPWR VPWR _1170_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload44 clknet_leaf_14_clk VGND VGND VPWR VPWR clkload44/Y sky130_fd_sc_hd__inv_6
Xclkload33 clknet_leaf_20_clk VGND VGND VPWR VPWR clkload33/X sky130_fd_sc_hd__clkbuf_1
Xclkload22 clknet_leaf_12_clk VGND VGND VPWR VPWR clkload22/Y sky130_fd_sc_hd__bufinv_16
X_6380_ clknet_leaf_81_clk _0187_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[4\] sky130_fd_sc_hd__dfrtp_1
X_3592_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1109_ sky130_fd_sc_hd__inv_2
X_5400_ tree_instances\[20\].u_tree.tree_state\[2\] tree_instances\[20\].u_tree.tree_state\[1\]
+ tree_instances\[20\].u_tree.tree_state\[0\] VGND VGND VPWR VPWR _2499_ sky130_fd_sc_hd__or3_1
Xclkload11 clknet_leaf_5_clk VGND VGND VPWR VPWR clkload11/Y sky130_fd_sc_hd__clkinvlp_4
X_5331_ _2438_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__clkbuf_1
Xclkload77 clknet_leaf_41_clk VGND VGND VPWR VPWR clkload77/Y sky130_fd_sc_hd__clkinv_2
Xclkload55 clknet_leaf_65_clk VGND VGND VPWR VPWR clkload55/Y sky130_fd_sc_hd__inv_6
Xclkload66 clknet_leaf_89_clk VGND VGND VPWR VPWR clkload66/Y sky130_fd_sc_hd__inv_6
XFILLER_0_11_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload88 clknet_leaf_51_clk VGND VGND VPWR VPWR clkload88/Y sky130_fd_sc_hd__bufinv_16
Xclkload99 clknet_leaf_63_clk VGND VGND VPWR VPWR clkload99/Y sky130_fd_sc_hd__clkinvlp_4
X_5262_ _2402_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__clkbuf_1
X_7001_ clknet_leaf_51_clk _0024_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5193_ tree_instances\[17\].u_tree.tree_state\[2\] tree_instances\[17\].u_tree.tree_state\[1\]
+ _2365_ VGND VGND VPWR VPWR _2366_ sky130_fd_sc_hd__or3_1
X_4213_ _1682_ _1671_ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__nor2_1
XANTENNA__6851__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4144_ _1617_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
X_4075_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1550_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_568 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_90_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_65_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6716_ clknet_leaf_46_clk _0464_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_18_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4977_ tree_instances\[13\].u_tree.frame_id_out\[4\] tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[13\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkload5 clknet_3_6__leaf_clk VGND VGND VPWR VPWR clkload5/Y sky130_fd_sc_hd__inv_2
X_3928_ _0758_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6647_ clknet_leaf_29_clk _0406_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3859_ _1341_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__clkbuf_1
X_6578_ clknet_leaf_49_clk _0347_ net35 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5529_ _2585_ VGND VGND VPWR VPWR _2586_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6939__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6521__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xload_slew28 net29 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_12
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_53_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_25_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5534__A0 _2589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6318__SET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6609__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_192 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5880_ _1227_ _2855_ _1820_ tree_instances\[1\].u_tree.ready_for_next VGND VGND VPWR
+ VPWR _0554_ sky130_fd_sc_hd__a22o_1
X_4900_ _1662_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[6\] _2179_
+ VGND VGND VPWR VPWR _2180_ sky130_fd_sc_hd__o21bai_1
Xclkbuf_leaf_72_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_4
X_4831_ tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[1\] _1830_ _0010_ VGND
+ VGND VPWR VPWR _2124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4762_ _2076_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3713_ _1212_ _1014_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__nor2_1
X_6501_ clknet_leaf_101_clk _0284_ net32 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4693_ _2033_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3644_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1154_ sky130_fd_sc_hd__clkbuf_1
X_6432_ clknet_leaf_98_clk _0225_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_31_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_43_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_95_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_101_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3575_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1093_ sky130_fd_sc_hd__buf_1
X_6363_ clknet_leaf_83_clk _0170_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_23_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5314_ tree_instances\[19\].u_tree.frame_id_out\[2\] tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _1252_ VGND VGND VPWR VPWR _2430_ sky130_fd_sc_hd__mux2_1
X_6294_ _0945_ _3101_ VGND VGND VPWR VPWR _3147_ sky130_fd_sc_hd__and2_1
X_5245_ _2393_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5750__A _2588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5176_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[6\] _2347_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ _1368_ _2349_ VGND VGND VPWR VPWR _2350_ sky130_fd_sc_hd__a221o_1
XANTENNA__4366__A _1112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4127_ _1585_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__clkbuf_1
X_4058_ _1531_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_39_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_63_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6773__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6702__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_54_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_435 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5507__B1 _0032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_194 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_107 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_438 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3360_ tree_instances\[19\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6443__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5030_ _2258_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3291_ _0835_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5570__A _2585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6981_ clknet_leaf_37_clk _0687_ net29 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5932_ _2916_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_0_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_0_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_45_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_64_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5863_ _2871_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4814_ _1276_ _2071_ VGND VGND VPWR VPWR _2115_ sky130_fd_sc_hd__and2_1
X_5794_ _2833_ _2443_ _2834_ VGND VGND VPWR VPWR _2835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4745_ tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[3\] _1835_ _0008_ VGND
+ VGND VPWR VPWR _2067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4676_ tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[2\] _1832_ _0006_ VGND
+ VGND VPWR VPWR _2023_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3627_ _0732_ tree_instances\[15\].u_tree.pipeline_valid\[0\] tree_instances\[15\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__o21a_1
X_6415_ clknet_leaf_2_clk _0216_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_31_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3558_ _1077_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6346_ clknet_leaf_20_clk _0153_ net26 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_8_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6277_ _3138_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__clkbuf_1
X_3489_ _1015_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__clkbuf_1
X_5228_ tree_instances\[17\].u_tree.frame_id_out\[1\] tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0909_ VGND VGND VPWR VPWR _2385_ sky130_fd_sc_hd__mux2_1
X_5159_ _0793_ VGND VGND VPWR VPWR _2333_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_36_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6954__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6652__SET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3175__A net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_27_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA__4779__B2 tree_instances\[11\].u_tree.ready_for_next VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_57_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_61_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_33_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6695__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_13_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5565__A _2588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6624__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4530_ _1934_ _1935_ _1937_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4461_ _0753_ _1884_ _0022_ tree_instances\[18\].u_tree.pipeline_valid\[0\] VGND
+ VGND VPWR VPWR _0128_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3412_ _0946_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6200_ _3095_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4392_ _1833_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_55 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6131_ _1327_ _2972_ VGND VGND VPWR VPWR _3047_ sky130_fd_sc_hd__and2_1
XFILLER_0_0_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3343_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _0884_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6062_ _2992_ _2995_ _3003_ _3004_ VGND VGND VPWR VPWR _3005_ sky130_fd_sc_hd__a31o_1
X_3274_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0821_ sky130_fd_sc_hd__clkbuf_1
X_5013_ tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[2\] _2125_ _0014_ VGND
+ VGND VPWR VPWR _2248_ sky130_fd_sc_hd__mux2_1
X_6964_ clknet_leaf_50_clk _0014_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_18_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_4
XPHY_EDGE_ROW_5_Right_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_101_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6895_ clknet_leaf_36_clk _0068_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5915_ _2157_ _2901_ VGND VGND VPWR VPWR _2908_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5846_ _1526_ _2427_ VGND VGND VPWR VPWR _2863_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5777_ _2447_ _2821_ _1020_ complete_votes\[0\] VGND VGND VPWR VPWR _2822_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__6365__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4728_ _2058_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4659_ _2014_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6329_ clknet_leaf_21_clk _0137_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_78_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_89_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3961_ _1061_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_18_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5700_ _2627_ _2739_ _2740_ _2744_ VGND VGND VPWR VPWR _2745_ sky130_fd_sc_hd__o211a_1
XFILLER_0_58_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3892_ _1219_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6805__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6680_ clknet_leaf_63_clk _0096_ net35 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
X_5631_ _2582_ tree_instances\[16\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2681_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_72_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5562_ _2585_ _2608_ _2609_ _2611_ tree_instances\[20\].u_tree.prediction_valid VGND
+ VGND VPWR VPWR _2612_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4513_ _1926_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_468 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5493_ _1197_ _1198_ _2550_ tree_instances\[20\].u_tree.ready_for_next VGND VGND
+ VPWR VPWR _0487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4444_ _1872_ _1851_ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_7_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4375_ _1821_ net17 VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__nor2_1
X_3326_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _0868_ sky130_fd_sc_hd__buf_1
XFILLER_0_95_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6114_ _3038_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6045_ _2949_ VGND VGND VPWR VPWR _2988_ sky130_fd_sc_hd__buf_1
X_3257_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[6\] tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[7\]
+ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__nand2_1
X_3188_ _0740_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5626__B_N _2578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6947_ clknet_leaf_88_clk _0659_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[0\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__6546__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6878_ clknet_leaf_12_clk _0597_ net29 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5829_ _2852_ VGND VGND VPWR VPWR _2853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6483__SET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_15_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_3_7__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_566 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4160_ _1116_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4091_ _1557_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6801_ clknet_leaf_43_clk _0523_ net36 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4993_ _2235_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__clkbuf_1
X_3944_ _1423_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__clkbuf_1
X_6732_ clknet_leaf_74_clk _0480_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.read_enable
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6663_ clknet_leaf_29_clk _0413_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_3875_ _1354_ _1358_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5614_ _2600_ tree_instances\[12\].u_tree.frame_id_out\[2\] _2662_ _2663_ tree_instances\[12\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2664_ sky130_fd_sc_hd__o221a_1
XFILLER_0_45_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6594_ clknet_leaf_60_clk _0358_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5545_ _2594_ _2596_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5476_ _0028_ VGND VGND VPWR VPWR _2550_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4427_ _1858_ _1851_ VGND VGND VPWR VPWR _1859_ sky130_fd_sc_hd__and2_1
X_4358_ _1803_ tree_instances\[8\].u_tree.pipeline_valid\[0\] tree_instances\[8\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__or3b_1
XFILLER_0_39_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4289_ _1756_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__clkbuf_1
X_3309_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _0852_ sky130_fd_sc_hd__buf_1
X_6028_ _2976_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6798__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_107_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6727__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6380__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_40_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5663__A _2631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_330 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_8_Left_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3627__A1 _0732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6468__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3660_ _1158_ _1161_ _1164_ _1168_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__or4_1
XFILLER_0_15_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload34 clknet_leaf_21_clk VGND VGND VPWR VPWR clkload34/Y sky130_fd_sc_hd__clkinv_1
XFILLER_0_70_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload12 clknet_leaf_6_clk VGND VGND VPWR VPWR clkload12/Y sky130_fd_sc_hd__inv_6
X_3591_ _1105_ _1107_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__nand2_1
Xclkload23 clknet_leaf_92_clk VGND VGND VPWR VPWR clkload23/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_35_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5330_ _1569_ _2414_ VGND VGND VPWR VPWR _2438_ sky130_fd_sc_hd__and2_1
Xclkload78 clknet_leaf_42_clk VGND VGND VPWR VPWR clkload78/Y sky130_fd_sc_hd__clkinv_4
Xclkload45 clknet_leaf_15_clk VGND VGND VPWR VPWR clkload45/Y sky130_fd_sc_hd__clkinv_2
Xclkload56 clknet_leaf_66_clk VGND VGND VPWR VPWR clkload56/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_2_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkload67 clknet_leaf_69_clk VGND VGND VPWR VPWR clkload67/Y sky130_fd_sc_hd__clkinv_1
XANTENNA__5573__A _2622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5261_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[2\] _1382_ _2399_
+ VGND VGND VPWR VPWR _2402_ sky130_fd_sc_hd__mux2_1
Xclkload89 clknet_leaf_52_clk VGND VGND VPWR VPWR clkload89/X sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_53_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5304__A1 _2249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_7000_ clknet_leaf_52_clk _0023_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4212_ _1677_ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__clkbuf_1
X_5192_ _0020_ VGND VGND VPWR VPWR _2365_ sky130_fd_sc_hd__inv_2
X_4143_ tree_instances\[0\].u_tree.prediction_valid _0737_ VGND VGND VPWR VPWR _1617_
+ sky130_fd_sc_hd__and2b_1
X_4074_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1549_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6891__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6820__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6715_ clknet_leaf_35_clk _0463_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_4976_ _2226_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3927_ _1406_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6646_ clknet_leaf_32_clk _0405_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkload6 clknet_3_7__leaf_clk VGND VGND VPWR VPWR clkload6/X sky130_fd_sc_hd__clkbuf_4
X_3858_ _1342_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6577_ clknet_leaf_49_clk _0346_ net35 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3789_ _1269_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5528_ current_voting_frame\[3\] VGND VGND VPWR VPWR _2585_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5459_ _1489_ _2534_ VGND VGND VPWR VPWR _2541_ sky130_fd_sc_hd__and2_1
XANTENNA__6979__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_70_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3178__A _0732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_376 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_519 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6649__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4830_ _2123_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4761_ tree_instances\[11\].u_tree.frame_id_out\[4\] tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[11\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3712_ _1013_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6500_ clknet_leaf_3_clk _0283_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.gen_tree_13.u_tree_rom.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_4692_ tree_instances\[10\].u_tree.frame_id_out\[2\] tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _1136_ VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__mux2_1
X_3643_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__clkbuf_1
X_6431_ clknet_leaf_100_clk _0224_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6362_ clknet_leaf_80_clk _0169_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5313_ _2429_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__clkbuf_1
X_3574_ _1091_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6293_ _3146_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__clkbuf_1
X_5244_ _1380_ _2314_ VGND VGND VPWR VPWR _2393_ sky130_fd_sc_hd__and2_1
X_5175_ _1371_ _2348_ VGND VGND VPWR VPWR _2349_ sky130_fd_sc_hd__nor2_1
X_4126_ _1574_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6319__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6890__SET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4057_ _1087_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_39_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_104_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5764__B2 _2589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5764__A1 _2619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6387__SET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_50_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4959_ _1837_ tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[4\] _1824_ VGND
+ VGND VPWR VPWR _2216_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_89_Left_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6629_ clknet_leaf_56_clk _0388_ net37 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6459__D _0034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_98_Left_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_119 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3290_ _0834_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND
+ VPWR VPWR _0835_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6412__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6980_ clknet_leaf_15_clk _0686_ net29 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5931_ tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[4\] tree_instances\[0\].u_tree.frame_id_in\[4\]
+ _0030_ VGND VGND VPWR VPWR _2916_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_0_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_36_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5862_ tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[4\] tree_instances\[0\].u_tree.frame_id_in\[4\]
+ _0026_ VGND VGND VPWR VPWR _2871_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_64_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4813_ _2114_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5746__A1 _2576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5793_ _2729_ _2820_ _2829_ complete_votes\[3\] _1018_ VGND VGND VPWR VPWR _2834_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_8_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4744_ _2066_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4675_ _2022_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__clkbuf_1
X_3626_ tree_instances\[15\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_341 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6414_ clknet_leaf_12_clk _0088_ net25 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
X_3557_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[4\] tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[5\]
+ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6345_ clknet_leaf_21_clk _0152_ net26 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_6276_ tree_instances\[6\].u_tree.frame_id_out\[4\] tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[6\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _3138_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_8_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3488_ _1013_ _1014_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__or2_1
X_5227_ _2384_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__clkbuf_1
X_5158_ _2331_ VGND VGND VPWR VPWR _2332_ sky130_fd_sc_hd__clkbuf_1
X_5089_ _2288_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__clkbuf_1
X_4109_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1584_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6748__SET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6994__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5671__A _2627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6923__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_load_slew33_A net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_33_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5728__B2 _2589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5728__A1 _2709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_61_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4460_ tree_instances\[18\].u_tree.tree_state\[0\] _0752_ VGND VGND VPWR VPWR _1884_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4391_ tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[2\] _1832_ _0040_ VGND
+ VGND VPWR VPWR _1833_ sky130_fd_sc_hd__mux2_1
X_3411_ _0944_ _0945_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3342_ _0866_ net17 tree_instances\[1\].u_tree.tree_state\[1\] VGND VGND VPWR VPWR
+ _0068_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6130_ _3046_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6061_ tree_instances\[5\].u_tree.read_enable VGND VGND VPWR VPWR _3004_ sky130_fd_sc_hd__inv_2
X_3273_ _0816_ _0819_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__nand2_1
X_5012_ _2247_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__clkbuf_1
X_6963_ clknet_leaf_49_clk _0013_ net35 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6894_ clknet_leaf_36_clk _0026_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5914_ _2907_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_101_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5845_ _2862_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5776_ _2729_ _2820_ VGND VGND VPWR VPWR _2821_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4727_ _1615_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[3\] _2010_
+ VGND VGND VPWR VPWR _2058_ sky130_fd_sc_hd__mux2_1
X_4658_ _1637_ _2012_ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3609_ _1122_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4589_ tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[0\] _1827_ _0044_ VGND
+ VGND VPWR VPWR _1969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6328_ clknet_leaf_22_clk _0136_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6334__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6259_ tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[2\] _2595_ _0038_ VGND
+ VGND VPWR VPWR _3129_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_11_Right_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_17_Left_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6135__B2 tree_instances\[4\].u_tree.ready_for_next VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_20_Right_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_26_Left_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3960_ _1435_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_18_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_35_Left_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_46_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3891_ _1360_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5576__A _2586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5630_ _2610_ tree_instances\[16\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2680_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_70_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6794__SET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5561_ _2610_ tree_instances\[20\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2611_
+ sky130_fd_sc_hd__xnor2_1
X_4512_ _1302_ _1839_ VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6845__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5492_ _2559_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_44_Left_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4443_ _1871_ VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4374_ _0865_ VGND VGND VPWR VPWR _1821_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3325_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _0867_ sky130_fd_sc_hd__buf_1
X_6113_ tree_instances\[4\].u_tree.frame_id_out\[2\] tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0849_ VGND VGND VPWR VPWR _3038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3256_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _0803_ sky130_fd_sc_hd__inv_2
X_6044_ _2985_ tree_instances\[3\].u_tree.node_data\[107\] _2987_ VGND VGND VPWR VPWR
+ _0611_ sky130_fd_sc_hd__a21o_1
X_3187_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[1\] tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[0\]
+ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__or2_1
XPHY_EDGE_ROW_53_Left_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6946_ clknet_leaf_25_clk _0658_ net24 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6877_ clknet_leaf_74_clk _0596_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_64_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5828_ _1932_ _1968_ VGND VGND VPWR VPWR _2852_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5759_ _2580_ _2801_ _2802_ _2803_ tree_instances\[6\].u_tree.prediction_valid VGND
+ VGND VPWR VPWR _2804_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_62_Left_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6586__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6515__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_73_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_71_Left_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_409 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5800__B1 _2583_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_43_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_283 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_80_Left_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_38 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_578 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4090_ _1559_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6800_ clknet_leaf_41_clk _0522_ net33 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4992_ _1684_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[3\] _2231_
+ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__mux2_1
X_6731_ clknet_leaf_35_clk _0479_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.current_node_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3943_ _1179_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6662_ clknet_leaf_33_clk _0412_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_3874_ _1356_ _1357_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_5613_ _2610_ tree_instances\[12\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2663_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6593_ clknet_leaf_59_clk _0357_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5544_ _2595_ _1834_ _2593_ VGND VGND VPWR VPWR _2596_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5475_ _0865_ VGND VGND VPWR VPWR _2549_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4426_ _0985_ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4530__B1 _1937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4357_ _1812_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__inv_2
X_4288_ _1747_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__clkbuf_1
X_3308_ _0850_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__clkbuf_1
X_3239_ _0784_ _0787_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__nand2_1
X_6027_ tree_instances\[3\].u_tree.frame_id_out\[3\] tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0799_ VGND VGND VPWR VPWR _2976_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_107_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6929_ clknet_leaf_16_clk _0102_ net29 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6767__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_40_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_20_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_526 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_109_Left_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6437__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload35 clknet_leaf_22_clk VGND VGND VPWR VPWR clkload35/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_70_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload13 clknet_leaf_7_clk VGND VGND VPWR VPWR clkload13/Y sky130_fd_sc_hd__clkinv_1
X_3590_ _1106_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__clkbuf_1
Xclkload24 clknet_leaf_93_clk VGND VGND VPWR VPWR clkload24/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_97_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload46 clknet_leaf_16_clk VGND VGND VPWR VPWR clkload46/Y sky130_fd_sc_hd__inv_6
Xclkload57 clknet_leaf_80_clk VGND VGND VPWR VPWR clkload57/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload68 clknet_leaf_70_clk VGND VGND VPWR VPWR clkload68/Y sky130_fd_sc_hd__clkinv_1
X_5260_ _2401_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__clkbuf_1
Xclkload79 clknet_leaf_43_clk VGND VGND VPWR VPWR clkload79/Y sky130_fd_sc_hd__inv_6
XFILLER_0_50_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4211_ _1680_ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__clkbuf_1
X_5191_ _2364_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4142_ _1616_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
X_4073_ _1548_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4975_ tree_instances\[13\].u_tree.frame_id_out\[3\] tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[3\]
+ tree_instances\[13\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6714_ clknet_leaf_34_clk _0462_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6860__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3926_ _1405_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6645_ clknet_leaf_34_clk _0404_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3857_ _1331_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__clkbuf_1
Xclkload7 clknet_leaf_0_clk VGND VGND VPWR VPWR clkload7/Y sky130_fd_sc_hd__inv_6
X_3788_ _1271_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6576_ clknet_leaf_61_clk _0345_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5527_ _2584_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__clkbuf_1
X_5458_ _2540_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__clkbuf_1
X_4409_ _1844_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
X_5389_ _2487_ VGND VGND VPWR VPWR _2491_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_70_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5059__A1 _2249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6948__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_25_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6530__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_81_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5298__A1 _2122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6689__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6618__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5222__A1 _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4760_ _2075_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3711_ _1210_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4691_ _2032_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__clkbuf_1
X_3642_ _1151_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6430_ clknet_leaf_97_clk _0223_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_70_278 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6361_ clknet_leaf_77_clk _0168_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_5312_ tree_instances\[19\].u_tree.frame_id_out\[1\] tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _1252_ VGND VGND VPWR VPWR _2429_ sky130_fd_sc_hd__mux2_1
X_3573_ tree_instances\[9\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_49_Right_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6292_ _2475_ _3101_ VGND VGND VPWR VPWR _3146_ sky130_fd_sc_hd__and2_1
X_5243_ _2392_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5174_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[2\] VGND VGND VPWR
+ VPWR _2348_ sky130_fd_sc_hd__inv_2
XANTENNA__6565__D _0040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4125_ _1594_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__clkbuf_1
X_4056_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1532_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_58_Right_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_104_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_50_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4958_ _2215_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__clkbuf_1
X_3909_ _1390_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_4889_ tree_instances\[13\].u_tree.u_tree_weight_rom.cache_valid VGND VGND VPWR VPWR
+ _2169_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6628_ clknet_leaf_57_clk _0387_ net37 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_67_Right_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_30_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_104_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6559_ clknet_leaf_4_clk _0333_ net26 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Right_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_58_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5669__A _2619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6782__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_52_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_85_Right_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_67_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_94_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_94_Right_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5691__A1 _2659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5930_ _2915_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6452__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_36_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5861_ _2870_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__clkbuf_1
X_4812_ _1275_ _2071_ VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__and2_1
X_5792_ _2443_ _1021_ VGND VGND VPWR VPWR _2833_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4743_ tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[2\] _1832_ _0008_ VGND
+ VGND VPWR VPWR _2066_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6413_ clknet_leaf_92_clk _0215_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
X_4674_ tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[1\] _1830_ _0006_ VGND
+ VGND VPWR VPWR _2022_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3625_ tree_instances\[10\].u_tree.tree_state\[0\] _1135_ _1136_ VGND VGND VPWR VPWR
+ _0047_ sky130_fd_sc_hd__a21o_1
X_3556_ _1075_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6344_ clknet_leaf_90_clk _0106_ net31 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
X_6275_ _3137_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__clkbuf_1
X_3487_ tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1014_ sky130_fd_sc_hd__buf_1
X_5226_ tree_instances\[17\].u_tree.frame_id_out\[0\] tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0909_ VGND VGND VPWR VPWR _2384_ sky130_fd_sc_hd__mux2_1
XANTENNA__5682__A1 _2583_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5157_ _2330_ VGND VGND VPWR VPWR _2331_ sky130_fd_sc_hd__clkbuf_1
X_5088_ _1083_ _2254_ VGND VGND VPWR VPWR _2288_ sky130_fd_sc_hd__and2_1
X_4108_ _1582_ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__clkbuf_1
X_4039_ _1515_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6963__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5673__A1 _2580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_175 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_33_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_61_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_13_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_245 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3410_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[8\] VGND VGND VPWR
+ VPWR _0945_ sky130_fd_sc_hd__clkbuf_1
X_4390_ tree_instances\[0\].u_tree.frame_id_in\[2\] VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__clkbuf_4
X_3341_ _0875_ _0882_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6060_ _1240_ _2996_ _2997_ _3000_ _3002_ VGND VGND VPWR VPWR _3003_ sky130_fd_sc_hd__o2111a_1
X_3272_ _0818_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND
+ VPWR VPWR _0819_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5011_ tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[1\] _2246_ _0014_ VGND
+ VGND VPWR VPWR _2247_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6633__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6962_ clknet_leaf_50_clk _0055_ net35 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_6893_ clknet_leaf_45_clk _0025_ net36 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5913_ _2160_ _2901_ VGND VGND VPWR VPWR _2907_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5844_ _1519_ _2427_ VGND VGND VPWR VPWR _2862_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_627 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5775_ _2764_ _2800_ _2819_ VGND VGND VPWR VPWR _2820_ sky130_fd_sc_hd__or3_2
XFILLER_0_44_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4726_ _2057_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4657_ _2013_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3608_ tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6327_ clknet_leaf_26_clk _0135_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4588_ _1917_ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__clkbuf_1
X_3539_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__clkbuf_1
X_6258_ _3128_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__clkbuf_1
X_6189_ _3080_ _3035_ VGND VGND VPWR VPWR _3090_ sky130_fd_sc_hd__and2_1
X_5209_ _2346_ _2367_ VGND VGND VPWR VPWR _2375_ sky130_fd_sc_hd__and2_1
XANTENNA__6374__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6303__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_67_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3467__A _0994_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_204 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_270 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_89_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkload0_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_18_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3890_ _1372_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5560_ current_voting_frame\[4\] VGND VGND VPWR VPWR _2610_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4511_ _1925_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5491_ tree_instances\[20\].u_tree.prediction_out tree_instances\[20\].u_tree.pipeline_prediction\[0\]\[0\]
+ tree_instances\[20\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4442_ _1870_ VGND VGND VPWR VPWR _1871_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6885__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4373_ _1820_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6814__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3324_ _0865_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__clkbuf_1
X_6112_ _3037_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__clkbuf_1
X_3255_ tree_instances\[2\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__clkbuf_1
X_6043_ tree_instances\[3\].u_tree.u_tree_weight_rom.gen_tree_3.u_tree_rom.node_data\[107\]
+ _2984_ _2986_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_data\[107\] VGND
+ VGND VPWR VPWR _2987_ sky130_fd_sc_hd__a22o_1
X_3186_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[3\] _0738_ VGND VGND
+ VPWR VPWR _0739_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6945_ clknet_leaf_26_clk _0657_ net24 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6876_ clknet_3_5__leaf_clk _0595_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5827_ _0737_ _2495_ _1818_ tree_instances\[0\].u_tree.ready_for_next VGND VGND VPWR
+ VPWR _0530_ sky130_fd_sc_hd__a22o_1
XFILLER_0_91_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5758_ _2622_ tree_instances\[6\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2803_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4709_ _1606_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[3\] tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ _1586_ _2043_ VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5689_ _2622_ _2732_ tree_instances\[9\].u_tree.frame_id_out\[4\] _2631_ _2733_ VGND
+ VGND VPWR VPWR _2734_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_73_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6555__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5628__A1 _2575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5677__A _2589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5800__A1 _2580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_15_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_43_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6522__SET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6585__SET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4991_ _2234_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5587__A _2585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6730_ clknet_leaf_68_clk _0478_ net36 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3942_ _1411_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6661_ clknet_leaf_34_clk _0411_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_3873_ _1219_ _1216_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_18_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6592_ clknet_leaf_34_clk _0356_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.cache_valid
+ sky130_fd_sc_hd__dfxtp_1
X_5612_ _2610_ tree_instances\[12\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2662_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_60_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5543_ tree_instances\[0\].u_tree.frame_id_in\[2\] VGND VGND VPWR VPWR _2595_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5526__S _1020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5474_ _2548_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5858__A1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4425_ _1857_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
X_4356_ _1803_ tree_instances\[7\].u_tree.pipeline_valid\[0\] tree_instances\[7\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1812_ sky130_fd_sc_hd__or3b_2
XFILLER_0_1_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3307_ tree_instances\[3\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__buf_1
X_4287_ _1754_ VGND VGND VPWR VPWR _1755_ sky130_fd_sc_hd__clkbuf_1
X_3238_ _0785_ _0786_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__nor2_1
X_6026_ _2975_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__clkbuf_1
X_3169_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _0725_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_93_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_107_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6928_ clknet_leaf_31_clk _0641_ net29 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XANTENNA__4597__A1 _1837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6859_ clknet_leaf_77_clk _0579_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_40_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6736__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_20_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_75_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_86_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_84_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_56_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload25 clknet_leaf_94_clk VGND VGND VPWR VPWR clkload25/Y sky130_fd_sc_hd__clkinv_1
Xclkload14 clknet_leaf_8_clk VGND VGND VPWR VPWR clkload14/Y sky130_fd_sc_hd__clkinvlp_2
Xclkload47 clknet_leaf_31_clk VGND VGND VPWR VPWR clkload47/Y sky130_fd_sc_hd__clkinv_2
Xclkload36 clknet_leaf_24_clk VGND VGND VPWR VPWR clkload36/Y sky130_fd_sc_hd__clkinv_1
Xclkload69 clknet_leaf_71_clk VGND VGND VPWR VPWR clkload69/Y sky130_fd_sc_hd__bufinv_16
XANTENNA__6477__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkload58 clknet_leaf_81_clk VGND VGND VPWR VPWR clkload58/Y sky130_fd_sc_hd__clkinv_2
XANTENNA__6406__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4210_ _1681_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__clkbuf_1
X_5190_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_data\[12\] tree_instances\[16\].u_tree.u_tree_weight_rom.gen_tree_16.u_tree_rom.node_data\[12\]
+ _2363_ VGND VGND VPWR VPWR _2364_ sky130_fd_sc_hd__mux2_1
X_4141_ tree_instances\[20\].u_tree.prediction_valid _1197_ VGND VGND VPWR VPWR _1616_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_48_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4072_ tree_instances\[19\].u_tree.prediction_valid _1252_ VGND VGND VPWR VPWR _1548_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_92_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4974_ _2225_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__clkbuf_1
X_6713_ clknet_leaf_47_clk _0461_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_86_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3925_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1405_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6644_ clknet_leaf_32_clk _0403_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload8 clknet_leaf_2_clk VGND VGND VPWR VPWR clkload8/Y sky130_fd_sc_hd__clkinv_4
X_3856_ _1334_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__clkbuf_1
X_3787_ _1268_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6575_ clknet_leaf_64_clk _0344_ net35 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5526_ _2583_ net4 _1020_ VGND VGND VPWR VPWR _2584_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5457_ _1480_ _2534_ VGND VGND VPWR VPWR _2540_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4408_ tree_instances\[7\].u_tree.frame_id_out\[3\] tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0970_ VGND VGND VPWR VPWR _1844_ sky130_fd_sc_hd__mux2_1
X_5388_ _2469_ VGND VGND VPWR VPWR _2490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_70_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4339_ _0730_ VGND VGND VPWR VPWR _1803_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6009_ _2964_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_66_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA__6008__A1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_25_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_53_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6988__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_81_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6917__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6570__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_57_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3710_ _1009_ _1209_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__nor2_1
XANTENNA__6658__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4690_ tree_instances\[10\].u_tree.frame_id_out\[1\] tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _1136_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__mux2_1
X_3641_ _1150_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3572_ _1080_ _1081_ _1085_ _1090_ tree_instances\[14\].u_tree.tree_state\[1\] VGND
+ VGND VPWR VPWR _0056_ sky130_fd_sc_hd__a41o_1
XFILLER_0_70_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6360_ clknet_leaf_81_clk _0167_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_87_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5311_ _2428_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6291_ _3145_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__clkbuf_1
X_5242_ _1384_ _2314_ VGND VGND VPWR VPWR _2392_ sky130_fd_sc_hd__and2_1
X_5173_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[6\] VGND VGND VPWR
+ VPWR _2347_ sky130_fd_sc_hd__inv_2
X_4124_ _1598_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__clkbuf_1
Xinput1 feature_valid VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_2
X_4055_ _1069_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_48_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_104_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_582 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6399__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4957_ _1835_ tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[3\] _1824_ VGND
+ VGND VPWR VPWR _2215_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3908_ tree_instances\[14\].u_tree.prediction_valid _0735_ VGND VGND VPWR VPWR _1390_
+ sky130_fd_sc_hd__and2b_1
X_4888_ _2168_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6328__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6627_ clknet_leaf_58_clk _0386_ net38 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3839_ _0852_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_30_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6558_ clknet_leaf_4_clk _0332_ net26 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5509_ _0755_ _2570_ _0030_ tree_instances\[2\].u_tree.pipeline_valid\[0\] VGND VGND
+ VPWR VPWR _0493_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6489_ clknet_leaf_3_clk _0272_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_prediction\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_58_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_39_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6751__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_94_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5860_ tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[3\] _1834_ _0026_ VGND
+ VGND VPWR VPWR _2870_ sky130_fd_sc_hd__mux2_1
XANTENNA__6839__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4811_ _2113_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5791_ state\[0\] _2447_ complete_votes\[3\] _2831_ _2832_ VGND VGND VPWR VPWR _0513_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_71_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4742_ _2065_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4673_ _2021_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3624_ tree_instances\[10\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__buf_2
X_6412_ clknet_leaf_93_clk _0214_ net25 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.prediction_out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3555_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[6\] tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[7\]
+ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5534__S _1020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6343_ clknet_leaf_86_clk _0151_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[8\].u_tree.ready_for_next sky130_fd_sc_hd__dfstp_1
X_3486_ tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1013_ sky130_fd_sc_hd__clkbuf_1
X_6274_ tree_instances\[6\].u_tree.frame_id_out\[3\] tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0932_ VGND VGND VPWR VPWR _3137_ sky130_fd_sc_hd__mux2_1
X_5225_ _2383_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5156_ _2329_ VGND VGND VPWR VPWR _2330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5087_ _2287_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__clkbuf_1
X_4107_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1582_ sky130_fd_sc_hd__clkbuf_1
X_4038_ _1513_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_644 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_614 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6509__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5989_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[1\] _1422_ _2899_
+ VGND VGND VPWR VPWR _2954_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_170 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_187 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_13_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3340_ _0876_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[6\] _0881_ VGND
+ VGND VPWR VPWR _0882_ sky130_fd_sc_hd__or3_1
X_5010_ _1829_ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__clkbuf_4
X_3271_ _0817_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6961_ clknet_leaf_35_clk _0672_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6673__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6892_ clknet_leaf_45_clk _0067_ net36 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_5912_ _2906_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__clkbuf_1
X_5843_ _2861_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6602__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_639 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5774_ _2687_ _2810_ _2817_ _2818_ VGND VGND VPWR VPWR _2819_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4725_ _1613_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[2\] _2010_
+ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4656_ _1627_ _2012_ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__and2_1
X_3607_ _1120_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__clkbuf_1
X_4587_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_data\[12\] _1966_ _1967_
+ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6326_ clknet_leaf_22_clk _0134_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3538_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1059_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3469_ tree_instances\[19\].u_tree.ready_for_next tree_instances\[18\].u_tree.ready_for_next
+ tree_instances\[20\].u_tree.ready_for_next _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__nand4_2
X_6257_ tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[1\] _1829_ _0038_ VGND
+ VGND VPWR VPWR _3128_ sky130_fd_sc_hd__mux2_1
X_6188_ _3089_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__clkbuf_1
X_5208_ _2374_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__clkbuf_1
X_5139_ tree_instances\[16\].u_tree.frame_id_out\[3\] tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _1023_ VGND VGND VPWR VPWR _2318_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_67_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_66_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3418__A1 _0733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5947__B _2553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_78_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_216 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_19_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_89_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_18_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4510_ _1313_ _1840_ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__and2_1
X_5490_ _2558_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4441_ _0972_ VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_53_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_9_Right_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4372_ _1112_ tree_instances\[1\].u_tree.pipeline_valid\[0\] tree_instances\[1\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1820_ sky130_fd_sc_hd__or3b_1
X_6111_ tree_instances\[4\].u_tree.frame_id_out\[1\] tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0849_ VGND VGND VPWR VPWR _3037_ sky130_fd_sc_hd__mux2_1
X_3323_ tree_instances\[1\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__buf_1
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_107_Right_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3254_ _0801_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
X_6042_ _2983_ VGND VGND VPWR VPWR _2986_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6854__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3185_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0738_ sky130_fd_sc_hd__clkbuf_1
X_6944_ clknet_leaf_26_clk _0656_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6875_ clknet_leaf_76_clk _0594_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_48_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5826_ _2851_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5757_ _2622_ tree_instances\[6\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2802_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_17_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4708_ _1581_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[1\] _1996_
+ _1157_ VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__o22a_1
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6833__SET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5688_ _2582_ tree_instances\[9\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2733_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_102_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4639_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[5\] tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__xor2_1
XFILLER_0_8_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6309_ clknet_leaf_29_clk _0118_ net28 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_73_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6595__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6524__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_15_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_43_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4990_ _1686_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[2\] _2231_
+ VGND VGND VPWR VPWR _2234_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3941_ _1420_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3872_ _1355_ _0926_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6660_ clknet_leaf_2_clk _0054_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6591_ clknet_leaf_37_clk _0355_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_prediction\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5611_ _2631_ tree_instances\[8\].u_tree.frame_id_out\[4\] _2655_ _2658_ _2660_ VGND
+ VGND VPWR VPWR _2661_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__5807__S _0004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5542_ _1832_ _2593_ _1835_ VGND VGND VPWR VPWR _2594_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_26_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5473_ tree_instances\[1\].u_tree.current_node_data\[12\] tree_instances\[1\].u_tree.node_data\[12\]
+ _0866_ VGND VGND VPWR VPWR _2548_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4424_ _1856_ _1851_ VGND VGND VPWR VPWR _1857_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4355_ _1811_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3306_ tree_instances\[4\].u_tree.tree_state\[0\] _0848_ _0849_ VGND VGND VPWR VPWR
+ _0075_ sky130_fd_sc_hd__a21o_1
X_4286_ _1753_ VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__clkbuf_1
X_3237_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _0786_ sky130_fd_sc_hd__clkbuf_1
X_6025_ tree_instances\[3\].u_tree.frame_id_out\[2\] tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0799_ VGND VGND VPWR VPWR _2975_ sky130_fd_sc_hd__mux2_1
X_3168_ _0723_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6927_ clknet_leaf_71_clk _0640_ net38 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6858_ clknet_leaf_78_clk _0578_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5809_ tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[1\] _2246_ _0004_ VGND
+ VGND VPWR VPWR _2843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_609 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6789_ clknet_leaf_69_clk _0070_ net38 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_75_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5724__A1_N _2603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5018__A tree_instances\[0\].u_tree.frame_id_in\[4\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_32_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6776__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6705__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_86_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5688__A _2582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_56_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_560 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload26 clknet_leaf_95_clk VGND VGND VPWR VPWR clkload26/Y sky130_fd_sc_hd__clkinvlp_4
Xclkload15 clknet_leaf_99_clk VGND VGND VPWR VPWR clkload15/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkload48 clknet_leaf_32_clk VGND VGND VPWR VPWR clkload48/Y sky130_fd_sc_hd__clkinv_4
XTAP_TAPCELL_ROW_97_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload37 clknet_leaf_25_clk VGND VGND VPWR VPWR clkload37/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_50_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload59 clknet_leaf_82_clk VGND VGND VPWR VPWR clkload59/Y sky130_fd_sc_hd__inv_6
XFILLER_0_23_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6446__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4140_ _1593_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__clkbuf_1
X_4071_ _1545_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4973_ tree_instances\[13\].u_tree.frame_id_out\[2\] tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _1114_ VGND VGND VPWR VPWR _2225_ sky130_fd_sc_hd__mux2_1
X_6712_ clknet_leaf_34_clk _0460_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3924_ _1397_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__clkbuf_1
X_6643_ clknet_leaf_33_clk _0402_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_500 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload9 clknet_leaf_3_clk VGND VGND VPWR VPWR clkload9/Y sky130_fd_sc_hd__clkinv_4
X_3855_ _1339_ _1336_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__nand2_1
X_3786_ _1266_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__clkbuf_1
X_6574_ clknet_leaf_65_clk _0343_ net35 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5525_ _2582_ VGND VGND VPWR VPWR _2583_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5456_ _2539_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4407_ _1843_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5700__A1 _2627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5387_ _2464_ _1247_ VGND VGND VPWR VPWR _2489_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_70_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4338_ _1802_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__buf_2
X_4269_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1737_ sky130_fd_sc_hd__clkbuf_1
X_6008_ tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[2\] _2595_ _0032_ VGND
+ VGND VPWR VPWR _2964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_325 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5767__A1 _2709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_59_Left_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_53_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5955__B _2553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xrst_buf rst_n VGND VGND VPWR VPWR tree_instances\[0\].u_tree.rst_n sky130_fd_sc_hd__buf_12
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6957__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_68_Left_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_211 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3640_ _1149_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND
+ VPWR VPWR _1150_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3571_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6698__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5310_ tree_instances\[19\].u_tree.frame_id_out\[0\] tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _1252_ VGND VGND VPWR VPWR _2428_ sky130_fd_sc_hd__mux2_1
XANTENNA__6627__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6290_ _2474_ _3102_ VGND VGND VPWR VPWR _3145_ sky130_fd_sc_hd__and2_1
XFILLER_0_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5241_ _2391_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_3_0__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5172_ _2345_ VGND VGND VPWR VPWR _2346_ sky130_fd_sc_hd__clkbuf_1
X_4123_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1598_ sky130_fd_sc_hd__inv_2
X_4054_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1530_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_50_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4956_ _2214_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__clkbuf_1
X_3907_ _1389_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4887_ _2165_ tree_instances\[13\].u_tree.pipeline_prediction\[0\]\[0\] _2167_ VGND
+ VGND VPWR VPWR _2168_ sky130_fd_sc_hd__mux2_1
X_6626_ clknet_leaf_59_clk _0385_ net38 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3838_ _0858_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__buf_1
XFILLER_0_61_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6557_ clknet_leaf_0_clk _0331_ net32 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6368__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3769_ _1259_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_5508_ tree_instances\[2\].u_tree.tree_state\[0\] _0754_ VGND VGND VPWR VPWR _2570_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6488_ clknet_leaf_94_clk _0078_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5439_ _2518_ VGND VGND VPWR VPWR _2528_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6098__S _0034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_58_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_2_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6791__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6720__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4810_ tree_instances\[12\].u_tree.u_tree_weight_rom.cache_valid _2112_ VGND VGND
+ VPWR VPWR _2113_ sky130_fd_sc_hd__or2_1
XFILLER_0_68_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5790_ _2820_ _2830_ _2447_ VGND VGND VPWR VPWR _2832_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4741_ tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[1\] _1830_ _0008_ VGND
+ VGND VPWR VPWR _2065_ sky130_fd_sc_hd__mux2_1
XANTENNA__6879__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4672_ tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[0\] _1827_ _0006_ VGND
+ VGND VPWR VPWR _2021_ sky130_fd_sc_hd__mux2_1
X_3623_ _0731_ tree_instances\[10\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _1135_ sky130_fd_sc_hd__or2_1
X_6411_ clknet_leaf_91_clk _0213_ net25 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5815__S _0004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6461__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3554_ _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6342_ clknet_leaf_93_clk _0150_ net27 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.prediction_out
+ sky130_fd_sc_hd__dfrtp_1
X_6273_ _3136_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__clkbuf_1
X_3485_ _1011_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__clkbuf_1
X_5224_ tree_instances\[16\].u_tree.current_node_data\[12\] tree_instances\[16\].u_tree.node_data\[12\]
+ _0912_ VGND VGND VPWR VPWR _2383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5155_ _2323_ VGND VGND VPWR VPWR _2329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5086_ _1082_ _2255_ VGND VGND VPWR VPWR _2287_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4106_ _1580_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__clkbuf_1
X_4037_ _1506_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_35_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5988_ _2953_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4939_ _1723_ _2133_ VGND VGND VPWR VPWR _2206_ sky130_fd_sc_hd__and2_1
XANTENNA__6549__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6609_ clknet_leaf_39_clk _0373_ net30 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_7_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5696__A _2582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_199 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_13_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3372__A1 _0732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3270_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _0817_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6960_ clknet_leaf_67_clk _0103_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[5\].u_tree.prediction_valid sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5911_ _2162_ _2901_ VGND VGND VPWR VPWR _2906_ sky130_fd_sc_hd__and2_1
X_6891_ clknet_leaf_13_clk _0101_ net30 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
X_5842_ _1516_ _2427_ VGND VGND VPWR VPWR _2861_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_32_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5773_ _2654_ net19 _2671_ _2645_ VGND VGND VPWR VPWR _2818_ sky130_fd_sc_hd__a211o_1
XANTENNA__6642__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4724_ _2056_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4655_ _2011_ VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_44_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3606_ _1116_ _1119_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_431 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4586_ _1902_ tree_instances\[8\].u_tree.u_tree_weight_rom.gen_tree_8.u_tree_rom.node_data\[12\]
+ _1918_ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__and3_1
X_6325_ clknet_leaf_22_clk _0133_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3537_ _1053_ _1057_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6256_ _3127_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__clkbuf_1
X_3468_ tree_instances\[15\].u_tree.ready_for_next tree_instances\[14\].u_tree.ready_for_next
+ tree_instances\[17\].u_tree.ready_for_next tree_instances\[16\].u_tree.ready_for_next
+ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__and4_1
X_6187_ _2565_ _3035_ VGND VGND VPWR VPWR _3089_ sky130_fd_sc_hd__and2_1
X_5207_ _2344_ _2367_ VGND VGND VPWR VPWR _2374_ sky130_fd_sc_hd__and2_1
X_3399_ _0933_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__clkbuf_1
X_5138_ _2317_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_67_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5069_ _2278_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6383__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6312__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_78_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_10_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_load_slew31_A tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_18_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_46_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4440_ _1869_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6110_ _3036_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4371_ _1819_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__inv_2
X_3322_ _0851_ _0854_ _0861_ _0864_ tree_instances\[3\].u_tree.tree_state\[1\] VGND
+ VGND VPWR VPWR _0074_ sky130_fd_sc_hd__a41o_1
X_3253_ _0799_ _0800_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__or2b_1
XPHY_EDGE_ROW_13_Left_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6041_ _2969_ VGND VGND VPWR VPWR _2985_ sky130_fd_sc_hd__clkbuf_1
X_3184_ tree_instances\[0\].u_tree.tree_state\[0\] _0736_ _0737_ VGND VGND VPWR VPWR
+ _0045_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_109_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6943_ clknet_leaf_25_clk _0655_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6894__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6823__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6874_ clknet_leaf_76_clk _0593_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_5825_ tree_instances\[0\].u_tree.frame_id_out\[4\] tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[0\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2851_ sky130_fd_sc_hd__mux2_1
XPHY_EDGE_ROW_22_Left_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5756_ tree_instances\[6\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2801_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5687_ tree_instances\[9\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2732_ sky130_fd_sc_hd__inv_2
X_4707_ _1609_ _1999_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ _1596_ _2004_ VGND VGND VPWR VPWR _2042_ sky130_fd_sc_hd__o221a_1
X_4638_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[7\] VGND VGND VPWR
+ VPWR _1996_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4569_ _1781_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[0\] _1957_
+ VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6308_ clknet_leaf_18_clk _0117_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_31_Left_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_73_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6239_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[2\] _2481_ _3116_
+ VGND VGND VPWR VPWR _3119_ sky130_fd_sc_hd__mux2_1
XANTENNA__4836__A1 _1835_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6564__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_40_Left_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_15_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_43_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5013__A1 _2125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3940_ _1176_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__clkbuf_1
X_3871_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1355_ sky130_fd_sc_hd__inv_2
XANTENNA_clkbuf_leaf_50_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6590_ clknet_leaf_84_clk _0084_ net31 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5610_ _2659_ tree_instances\[8\].u_tree.frame_id_out\[3\] tree_instances\[8\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2660_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5541_ _1832_ _2593_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_65_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5472_ _2547_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__clkbuf_1
X_4423_ _1855_ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4354_ _1803_ tree_instances\[6\].u_tree.pipeline_valid\[0\] tree_instances\[6\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__or3b_1
XFILLER_0_22_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3305_ tree_instances\[4\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__buf_2
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4285_ _1093_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__clkbuf_1
X_6024_ _2974_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__clkbuf_1
X_3236_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _0785_ sky130_fd_sc_hd__clkbuf_1
X_3167_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _0723_ sky130_fd_sc_hd__clkbuf_1
X_6926_ clknet_leaf_72_clk _0639_ net38 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_18_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6857_ clknet_leaf_79_clk _0577_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5808_ _2842_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6788_ clknet_leaf_69_clk _0028_ net38 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5739_ _2579_ tree_instances\[14\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2784_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_364 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_481 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_75_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_20_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6745__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_86_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_86_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload16 clknet_leaf_100_clk VGND VGND VPWR VPWR clkload16/Y sky130_fd_sc_hd__clkinv_2
Xclkload49 clknet_leaf_33_clk VGND VGND VPWR VPWR clkload49/Y sky130_fd_sc_hd__inv_6
XFILLER_0_106_572 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload38 clknet_leaf_26_clk VGND VGND VPWR VPWR clkload38/Y sky130_fd_sc_hd__clkinv_1
Xclkload27 clknet_leaf_96_clk VGND VGND VPWR VPWR clkload27/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_206 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4070_ _1537_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6486__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6415__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4972_ _2224_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__clkbuf_1
X_6711_ clknet_leaf_48_clk _0459_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3923_ _1402_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6642_ clknet_leaf_34_clk _0401_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3854_ _1187_ _1323_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3785_ _1261_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__clkbuf_1
X_6573_ clknet_leaf_65_clk _0342_ net36 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5524_ current_voting_frame\[2\] VGND VGND VPWR VPWR _2582_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5455_ _1495_ _2534_ VGND VGND VPWR VPWR _2539_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4406_ tree_instances\[7\].u_tree.frame_id_out\[2\] tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0970_ VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5386_ _2470_ _2454_ VGND VGND VPWR VPWR _2488_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_70_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4337_ tree_instances\[20\].u_tree.pipeline_valid\[0\] tree_instances\[20\].u_tree.tree_state\[0\]
+ net1 VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__and3b_1
X_4268_ _1735_ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__clkbuf_1
X_3219_ _0768_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__clkbuf_1
X_6007_ _2963_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__clkbuf_1
X_4199_ _1670_ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5216__A1 _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_25_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6909_ clknet_leaf_37_clk _0622_ net29 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6926__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_5_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_587 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3570_ _1088_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_142 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5240_ _1382_ _2314_ VGND VGND VPWR VPWR _2391_ sky130_fd_sc_hd__and2_1
XANTENNA__5143__A0 tree_instances\[16\].u_tree.prediction_out VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_87_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5171_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _2345_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_18_Right_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4122_ _1162_ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__clkbuf_1
X_4053_ _1070_ VGND VGND VPWR VPWR _1529_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_27_Right_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4957__A0 _1835_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4955_ _1832_ tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[2\] _1824_ VGND
+ VGND VPWR VPWR _2214_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_50_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3906_ tree_instances\[13\].u_tree.prediction_valid _1114_ VGND VGND VPWR VPWR _1389_
+ sky130_fd_sc_hd__and2b_1
X_4886_ tree_instances\[13\].u_tree.tree_state\[0\] _1113_ _2166_ _0011_ VGND VGND
+ VPWR VPWR _2167_ sky130_fd_sc_hd__a211o_1
XFILLER_0_46_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6625_ clknet_leaf_58_clk _0384_ net38 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3837_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1322_ sky130_fd_sc_hd__inv_2
X_3768_ tree_instances\[7\].u_tree.prediction_valid _0970_ VGND VGND VPWR VPWR _1259_
+ sky130_fd_sc_hd__and2b_1
X_6556_ clknet_leaf_0_clk _0330_ net32 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5507_ _0799_ _0800_ _0032_ tree_instances\[3\].u_tree.pipeline_valid\[0\] VGND VGND
+ VPWR VPWR _0492_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3699_ _1149_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5634__A_N _2578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_5_Left_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6487_ clknet_leaf_87_clk _0036_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5438_ _2527_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_36_Right_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5369_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _2471_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6337__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_315 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_38_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_45_Right_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_54_Right_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6760__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_63_Right_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4740_ _2064_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4671_ _2020_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3622_ _1121_ _1134_ _1115_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_71_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6410_ clknet_leaf_91_clk _0212_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_72_Right_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6341_ clknet_leaf_94_clk _0149_ net31 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3553_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[1\] tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[2\]
+ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__or2_1
XANTENNA__6848__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3484_ _1010_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__clkbuf_1
X_6272_ tree_instances\[6\].u_tree.frame_id_out\[2\] tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0932_ VGND VGND VPWR VPWR _3136_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5223_ _2382_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__clkbuf_1
X_5154_ _2327_ VGND VGND VPWR VPWR _2328_ sky130_fd_sc_hd__clkbuf_1
X_4105_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1580_ sky130_fd_sc_hd__inv_2
X_5085_ _2286_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_87_Left_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_81_Right_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4036_ _0891_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5987_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[0\] _1407_ _2899_
+ VGND VGND VPWR VPWR _2953_ sky130_fd_sc_hd__mux2_1
X_4938_ _2205_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4869_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _2150_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_90_Right_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6608_ clknet_leaf_39_clk _0372_ net30 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_462 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6589__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6539_ clknet_leaf_4_clk _0313_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_30_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6518__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_7_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xmax_cap21 _2577_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_97_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3497__A _0732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_510 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6941__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5910_ _2905_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_49_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6890_ clknet_leaf_71_clk _0609_ net36 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
X_5841_ _2860_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4388__A1 _1830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_60_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5772_ _2812_ _2816_ _2624_ _2613_ VGND VGND VPWR VPWR _2817_ sky130_fd_sc_hd__a211o_1
XFILLER_0_8_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_32_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3200__A _0733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4723_ _1607_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[1\] _2010_
+ VGND VGND VPWR VPWR _2056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4654_ tree_instances\[0\].u_tree.tree_state\[1\] tree_instances\[0\].u_tree.tree_state\[2\]
+ _1818_ VGND VGND VPWR VPWR _2011_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3605_ _1118_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6682__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4585_ _1957_ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6611__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6324_ clknet_leaf_23_clk _0132_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3536_ _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6255_ tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[0\] _1826_ _0038_ VGND
+ VGND VPWR VPWR _3127_ sky130_fd_sc_hd__mux2_1
X_5206_ _2373_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__clkbuf_1
X_3467_ _0994_ _0995_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6186_ _3088_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_95_Left_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3398_ tree_instances\[5\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__buf_1
X_5137_ tree_instances\[16\].u_tree.frame_id_out\[2\] tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _1023_ VGND VGND VPWR VPWR _2317_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5068_ tree_instances\[15\].u_tree.frame_id_out\[2\] tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _1137_ VGND VGND VPWR VPWR _2278_ sky130_fd_sc_hd__mux2_1
X_4019_ _1493_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_67_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_0_Right_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_78_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6352__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5554__A1_N _2600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_89_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_18_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_46_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5507__A1_N _0799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_354 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4370_ _1112_ tree_instances\[10\].u_tree.pipeline_valid\[0\] tree_instances\[10\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__or3b_1
XFILLER_0_110_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3321_ _0863_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3252_ _0732_ tree_instances\[3\].u_tree.pipeline_valid\[0\] tree_instances\[3\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6040_ _2949_ VGND VGND VPWR VPWR _2984_ sky130_fd_sc_hd__clkbuf_1
X_3183_ tree_instances\[0\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__buf_2
XFILLER_0_28_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_109_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6942_ clknet_leaf_26_clk _0654_ net24 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6873_ clknet_leaf_78_clk _0592_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_76_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5824_ _2850_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5755_ _2766_ _2771_ _2780_ _2799_ VGND VGND VPWR VPWR _2800_ sky130_fd_sc_hd__o211ai_2
XANTENNA__6863__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5686_ _2713_ tree_instances\[9\].u_tree.frame_id_out\[1\] tree_instances\[9\].u_tree.frame_id_out\[4\]
+ _2708_ VGND VGND VPWR VPWR _2731_ sky130_fd_sc_hd__o22a_1
X_4706_ _2037_ _2038_ _2039_ _2040_ _1997_ VGND VGND VPWR VPWR _2041_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4637_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[1\] VGND VGND VPWR
+ VPWR _1995_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4568_ _1956_ VGND VGND VPWR VPWR _1957_ sky130_fd_sc_hd__buf_1
XFILLER_0_40_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4499_ _1919_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
X_6307_ clknet_leaf_40_clk _0116_ net30 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3519_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1041_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_73_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6238_ _3118_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__clkbuf_1
X_6169_ _2567_ VGND VGND VPWR VPWR _3077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_96_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_15_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_43_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_87_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_4
X_3870_ _1353_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6201__A1 _1829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5540_ _2592_ _2593_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_11_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5471_ tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[4\] _2251_ _0028_ VGND
+ VGND VPWR VPWR _2547_ sky130_fd_sc_hd__mux2_1
X_4422_ _1854_ VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4353_ _1810_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__inv_2
X_3304_ _0733_ tree_instances\[4\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _0848_ sky130_fd_sc_hd__or2_1
X_4284_ _1751_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__clkbuf_1
X_3235_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__clkbuf_1
X_6023_ tree_instances\[3\].u_tree.frame_id_out\[1\] tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0799_ VGND VGND VPWR VPWR _2974_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_78_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_4
X_3166_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[8\] VGND VGND VPWR
+ VPWR _0722_ sky130_fd_sc_hd__inv_2
X_6925_ clknet_leaf_72_clk _0638_ net39 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6856_ clknet_leaf_66_clk _0576_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[2\].u_tree.frame_id_out\[4\] sky130_fd_sc_hd__dfrtp_1
X_3999_ _0879_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__clkbuf_1
X_5807_ tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[0\] _1826_ _0004_ VGND
+ VGND VPWR VPWR _2842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6787_ clknet_leaf_69_clk _0027_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5738_ tree_instances\[14\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2783_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_493 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_20_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5669_ _2619_ VGND VGND VPWR VPWR _2714_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_75_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_102_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6259__A1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_69_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_86_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6785__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4745__A1 _1835_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkload17 clknet_leaf_101_clk VGND VGND VPWR VPWR clkload17/Y sky130_fd_sc_hd__clkinvlp_4
XFILLER_0_106_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkload39 clknet_leaf_27_clk VGND VGND VPWR VPWR clkload39/Y sky130_fd_sc_hd__clkinv_2
XTAP_TAPCELL_ROW_97_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkload28 clknet_leaf_97_clk VGND VGND VPWR VPWR clkload28/Y sky130_fd_sc_hd__clkinv_4
XFILLER_0_2_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_0_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_106_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4971_ tree_instances\[13\].u_tree.frame_id_out\[1\] tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _1114_ VGND VGND VPWR VPWR _2224_ sky130_fd_sc_hd__mux2_1
X_6710_ clknet_leaf_47_clk _0458_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6455__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3922_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1402_ sky130_fd_sc_hd__inv_2
XFILLER_0_86_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6641_ clknet_leaf_62_clk _0400_ net37 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3853_ _1332_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3784_ _1273_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__clkbuf_1
X_6572_ clknet_leaf_65_clk _0341_ net35 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5523_ _2581_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5454_ _2538_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4405_ _1842_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5385_ _2455_ _2462_ VGND VGND VPWR VPWR _2487_ sky130_fd_sc_hd__nor2_1
X_4336_ _1801_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_70_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4267_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1735_ sky130_fd_sc_hd__clkbuf_1
X_3218_ _0765_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__or2_1
X_4198_ _1657_ _1665_ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__nand2_1
X_6006_ tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[1\] _1829_ _0032_ VGND
+ VGND VPWR VPWR _2963_ sky130_fd_sc_hd__mux2_1
X_3149_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _0705_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_53_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6908_ clknet_leaf_70_clk _0621_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.cached_data\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6839_ clknet_leaf_86_clk _0559_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_81_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_92_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_5_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_64_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_79_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_599 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_66 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5170_ _2343_ VGND VGND VPWR VPWR _2344_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4121_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1596_ sky130_fd_sc_hd__inv_2
X_4052_ _1528_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6636__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3203__A _0733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5705__A2_N _2606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4954_ _2213_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_1
X_3905_ _1387_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4885_ tree_instances\[13\].u_tree.tree_state\[1\] _0967_ tree_instances\[13\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _2166_ sky130_fd_sc_hd__nor3_1
X_6624_ clknet_leaf_57_clk _0383_ net37 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3836_ _1318_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__clkbuf_1
X_3767_ _0751_ _1254_ _1258_ tree_instances\[18\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0064_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6555_ clknet_leaf_1_clk _0329_ net26 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5506_ tree_instances\[11\].u_tree.tree_state\[0\] _0951_ _2569_ tree_instances\[11\].u_tree.pipeline_valid\[0\]
+ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__o22a_1
XTAP_TAPCELL_ROW_30_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3698_ _1143_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6486_ clknet_leaf_83_clk _0035_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5437_ _1498_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[7\] _2518_
+ VGND VGND VPWR VPWR _2527_ sky130_fd_sc_hd__mux2_1
X_5368_ _0937_ VGND VGND VPWR VPWR _2470_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5299_ _2421_ VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4319_ _1785_ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_58_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6377__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6306__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_38_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_106_Left_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_38_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5125__A1 _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_103_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4670_ _1634_ _2011_ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_363 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3621_ _1115_ _1121_ _1134_ tree_instances\[0\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0046_ sky130_fd_sc_hd__a31o_1
X_3552_ _1071_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_58 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6340_ clknet_leaf_90_clk _0148_ net31 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3483_ _1009_ tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND
+ VPWR VPWR _1010_ sky130_fd_sc_hd__or2_1
X_6271_ _3135_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__clkbuf_1
X_5222_ tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[4\] _2251_ _0020_ VGND
+ VGND VPWR VPWR _2382_ sky130_fd_sc_hd__mux2_1
XANTENNA__6888__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6817__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5153_ _0781_ VGND VGND VPWR VPWR _2327_ sky130_fd_sc_hd__clkbuf_1
X_4104_ _1578_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__clkbuf_1
X_5084_ _1543_ _2255_ VGND VGND VPWR VPWR _2286_ sky130_fd_sc_hd__and2_1
XANTENNA__6470__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4035_ _1505_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_360 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_35_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5986_ _2952_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4937_ _1713_ _2133_ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4868_ _2145_ VGND VGND VPWR VPWR _2149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6607_ clknet_leaf_37_clk _0371_ net30 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3819_ _1307_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4799_ _0839_ _2091_ VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6538_ clknet_leaf_4_clk _0312_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_6469_ clknet_leaf_28_clk _0257_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_7_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6558__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_102_Right_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6981__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6910__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6299__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5840_ _1512_ _2427_ VGND VGND VPWR VPWR _2860_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_511 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5771_ _2713_ tree_instances\[7\].u_tree.frame_id_out\[1\] _2814_ _2815_ tree_instances\[7\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2816_ sky130_fd_sc_hd__o2111a_1
XTAP_TAPCELL_ROW_60_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5585__A1 _2589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_32_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4722_ _2055_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4653_ _1994_ _2010_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__nand2_1
X_3604_ tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[6\] _1117_ VGND VGND
+ VPWR VPWR _1118_ sky130_fd_sc_hd__or2_1
X_4584_ _1965_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
X_6323_ clknet_leaf_22_clk _0131_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3535_ _1055_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3466_ tree_instances\[7\].u_tree.ready_for_next tree_instances\[6\].u_tree.ready_for_next
+ tree_instances\[9\].u_tree.ready_for_next tree_instances\[8\].u_tree.ready_for_next
+ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6254_ _3126_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__clkbuf_1
X_5205_ _2340_ _2367_ VGND VGND VPWR VPWR _2373_ sky130_fd_sc_hd__and2_1
X_6185_ _1885_ _3035_ VGND VGND VPWR VPWR _3088_ sky130_fd_sc_hd__and2_1
X_3397_ tree_instances\[6\].u_tree.tree_state\[0\] _0931_ _0932_ VGND VGND VPWR VPWR
+ _0079_ sky130_fd_sc_hd__a21o_1
XANTENNA__6651__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5136_ _2316_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__clkbuf_1
X_5067_ _2277_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__clkbuf_1
X_4018_ _1482_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_67_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5969_ _2936_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_78_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5037__B _2222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6321__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_89_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_127 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4831__S _0010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3320_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[7\] _0862_ VGND VGND
+ VPWR VPWR _0863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6409__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3251_ tree_instances\[3\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__buf_2
XFILLER_0_28_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3182_ _0733_ tree_instances\[0\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _0736_ sky130_fd_sc_hd__or2_1
XFILLER_0_28_53 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6941_ clknet_leaf_27_clk _0653_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_109_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6872_ clknet_leaf_78_clk _0591_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5823_ tree_instances\[0\].u_tree.frame_id_out\[3\] tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0737_ VGND VGND VPWR VPWR _2850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4741__S _0008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5754_ _2781_ _2788_ _2798_ VGND VGND VPWR VPWR _2799_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5685_ tree_instances\[9\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2730_ sky130_fd_sc_hd__inv_2
X_4705_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[6\] tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ VGND VGND VPWR VPWR _2040_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4636_ tree_instances\[10\].u_tree.u_tree_weight_rom.cache_valid VGND VGND VPWR VPWR
+ _1994_ sky130_fd_sc_hd__inv_2
XANTENNA__6832__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5730__A1 _2576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5730__B2 _2588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6306_ clknet_leaf_40_clk _0115_ net30 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4567_ tree_instances\[8\].u_tree.read_enable _1917_ VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__nand2_4
X_4498_ _1290_ _1840_ VGND VGND VPWR VPWR _1919_ sky130_fd_sc_hd__and2_1
X_3518_ _1039_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND
+ VPWR VPWR _1040_ sky130_fd_sc_hd__or2_1
X_3449_ _0977_ _0978_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_73_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6237_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[1\] _2486_ _3116_
+ VGND VGND VPWR VPWR _3118_ sky130_fd_sc_hd__mux2_1
X_6168_ _3075_ VGND VGND VPWR VPWR _3076_ sky130_fd_sc_hd__clkbuf_1
X_5119_ tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[1\] _2246_ _0018_ VGND
+ VGND VPWR VPWR _2306_ sky130_fd_sc_hd__mux2_1
X_6099_ _3029_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_15_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5721__A1 _2708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6573__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6502__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5470_ _2546_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4421_ _1853_ VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4352_ _1803_ tree_instances\[12\].u_tree.pipeline_valid\[0\] tree_instances\[12\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__or3b_1
X_4283_ _1094_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__clkbuf_1
X_3303_ _0844_ _0847_ tree_instances\[12\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR
+ _0009_ sky130_fd_sc_hd__o21a_1
X_3234_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _0783_ sky130_fd_sc_hd__inv_2
X_6022_ _2973_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__clkbuf_1
X_3165_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6924_ clknet_leaf_72_clk _0637_ net39 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6855_ clknet_leaf_66_clk _0575_ net36 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3998_ _0877_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5806_ _2589_ _2839_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__xnor2_1
X_6786_ clknet_leaf_69_clk _0069_ net38 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_91_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5737_ tree_instances\[14\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2782_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5668_ _2603_ VGND VGND VPWR VPWR _2713_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_20_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5703__B2 _2659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5599_ tree_instances\[1\].u_tree.frame_id_out\[3\] _2585_ VGND VGND VPWR VPWR _2649_
+ sky130_fd_sc_hd__or2b_1
X_4619_ _1800_ _1937_ VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_56_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6754__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_97_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkload18 clknet_leaf_102_clk VGND VGND VPWR VPWR clkload18/Y sky130_fd_sc_hd__clkinv_4
Xclkload29 clknet_leaf_98_clk VGND VGND VPWR VPWR clkload29/X sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_106_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4970_ _2223_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3921_ _1183_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6640_ clknet_leaf_62_clk _0399_ net35 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3852_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[5\] tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[6\]
+ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__nor2_1
X_6571_ clknet_leaf_61_clk _0340_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3783_ _1272_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__clkbuf_1
X_5522_ _2580_ net3 _1020_ VGND VGND VPWR VPWR _2581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6424__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5453_ _1497_ _2534_ VGND VGND VPWR VPWR _2538_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4404_ tree_instances\[7\].u_tree.frame_id_out\[1\] tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0970_ VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5384_ _2471_ VGND VGND VPWR VPWR _2486_ sky130_fd_sc_hd__clkbuf_1
X_4335_ _0731_ tree_instances\[18\].u_tree.pipeline_valid\[0\] tree_instances\[18\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1801_ sky130_fd_sc_hd__or3b_1
XFILLER_0_5_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_70_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4266_ _1733_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6005_ _2962_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__clkbuf_1
X_3217_ _0766_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__clkbuf_1
X_4197_ _1668_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4672__A1 _1827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_19_Left_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6907_ clknet_leaf_61_clk _0620_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_53_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_81_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6838_ clknet_leaf_85_clk _0558_ net39 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6769_ clknet_leaf_11_clk _0503_ net29 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.frame_id_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_28_Left_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_185 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5045__B _2222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6935__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_228 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_78 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4120_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1595_ sky130_fd_sc_hd__inv_2
X_4051_ tree_instances\[18\].u_tree.prediction_valid _0753_ VGND VGND VPWR VPWR _1528_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_36_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5603__B1 _2652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6676__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4953_ _1830_ tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[1\] _1824_ VGND
+ VGND VPWR VPWR _2213_ sky130_fd_sc_hd__mux2_1
X_3904_ _0915_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6605__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_50_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6006__S _0032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6623_ clknet_leaf_57_clk _0382_ net37 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4884_ tree_instances\[13\].u_tree.tree_state\[1\] tree_instances\[13\].u_tree.current_node_data\[12\]
+ tree_instances\[13\].u_tree.node_data\[12\] _2164_ VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3835_ _1189_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__clkbuf_1
X_3766_ _1257_ _0744_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__nor2_1
X_6554_ clknet_leaf_0_clk _0328_ net32 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5505_ tree_instances\[11\].u_tree.tree_state\[3\] _1816_ VGND VGND VPWR VPWR _2569_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_30_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_604 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6485_ clknet_leaf_86_clk _0077_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_5436_ _2526_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__clkbuf_1
X_3697_ _1199_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
X_5367_ _2466_ VGND VGND VPWR VPWR _2469_ sky130_fd_sc_hd__clkbuf_1
X_5298_ tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[0\] _2122_ _0024_ VGND
+ VGND VPWR VPWR _2421_ sky130_fd_sc_hd__mux2_1
X_4318_ _1048_ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_58_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4249_ _1717_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_38_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6346__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_258 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_494 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3304__A _0733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4834__S _0010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5061__A1 _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3620_ _1124_ _1133_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3551_ _1069_ _1070_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_291 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3482_ tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1009_ sky130_fd_sc_hd__buf_1
X_6270_ tree_instances\[6\].u_tree.frame_id_out\[1\] tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0932_ VGND VGND VPWR VPWR _3135_ sky130_fd_sc_hd__mux2_1
X_5221_ _2381_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5152_ _0785_ VGND VGND VPWR VPWR _2326_ sky130_fd_sc_hd__clkbuf_1
X_4103_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1578_ sky130_fd_sc_hd__inv_2
X_5083_ _2285_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4034_ _1501_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6857__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_63_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_35_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5985_ tree_instances\[3\].u_tree.u_tree_weight_rom.cache_valid _2951_ VGND VGND
+ VPWR VPWR _2952_ sky130_fd_sc_hd__or2_1
X_4936_ _2204_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4867_ _2143_ VGND VGND VPWR VPWR _2148_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6606_ clknet_leaf_35_clk _0370_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.read_enable
+ sky130_fd_sc_hd__dfrtp_1
X_3818_ _1306_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_420 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4798_ _1711_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[4\] VGND
+ VGND VPWR VPWR _2101_ sky130_fd_sc_hd__or2_1
X_6537_ clknet_leaf_4_clk _0311_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_104_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3749_ _0937_ _0939_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__nor2_1
X_6468_ clknet_leaf_28_clk _0256_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_63_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5419_ _2512_ _2513_ _2515_ VGND VGND VPWR VPWR _2516_ sky130_fd_sc_hd__or3b_1
X_6399_ clknet_leaf_51_clk _0201_ net35 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_7_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_78_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6598__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6527__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_640 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_150 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_16_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4829__S _0010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6950__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5770_ _2598_ tree_instances\[7\].u_tree.frame_id_out\[0\] tree_instances\[7\].u_tree.frame_id_out\[1\]
+ _2603_ VGND VGND VPWR VPWR _2815_ sky130_fd_sc_hd__a22oi_1
XTAP_TAPCELL_ROW_60_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4721_ _1591_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[0\] _2010_
+ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4652_ _2009_ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3603_ tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1117_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4583_ _1784_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[7\] _1956_
+ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__mux2_1
X_3534_ _1054_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND
+ VPWR VPWR _1055_ sky130_fd_sc_hd__or2_1
X_6322_ clknet_leaf_78_clk _0130_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.cache_valid
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4739__S _0008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6253_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_data\[107\] tree_instances\[5\].u_tree.u_tree_weight_rom.gen_tree_5.u_tree_rom.node_data\[107\]
+ _3125_ VGND VGND VPWR VPWR _3126_ sky130_fd_sc_hd__mux2_1
X_3465_ tree_instances\[11\].u_tree.ready_for_next tree_instances\[10\].u_tree.ready_for_next
+ tree_instances\[13\].u_tree.ready_for_next tree_instances\[12\].u_tree.ready_for_next
+ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__and4_1
X_5204_ _2372_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6184_ _3087_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__clkbuf_1
X_3396_ tree_instances\[6\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__buf_2
X_5135_ tree_instances\[16\].u_tree.frame_id_out\[1\] tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _1023_ VGND VGND VPWR VPWR _2316_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6691__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5066_ tree_instances\[15\].u_tree.frame_id_out\[1\] tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _1137_ VGND VGND VPWR VPWR _2277_ sky130_fd_sc_hd__mux2_1
X_4017_ _1487_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5273__A1 _2122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6620__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5968_ tree_instances\[3\].u_tree.pipeline_prediction\[0\]\[0\] _2933_ _2935_ VGND
+ VGND VPWR VPWR _2936_ sky130_fd_sc_hd__mux2_1
X_4919_ _2195_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5899_ _2898_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_78_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6779__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4384__S _0040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5016__A1 _2249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_111_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _0776_ _0779_ _0798_ tree_instances\[17\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0062_ sky130_fd_sc_hd__a31o_1
X_3181_ tree_instances\[14\].u_tree.tree_state\[0\] _0734_ _0735_ VGND VGND VPWR VPWR
+ _0055_ sky130_fd_sc_hd__a21o_1
XANTENNA__6449__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6940_ clknet_leaf_27_clk _0652_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6613__SET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_109_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6871_ clknet_leaf_79_clk _0590_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_5822_ _2849_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_17_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5753_ _2791_ _2793_ _2797_ VGND VGND VPWR VPWR _2798_ sky130_fd_sc_hd__and3_1
XFILLER_0_56_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4704_ _1573_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[6\] VGND
+ VGND VPWR VPWR _2039_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5684_ net10 VGND VGND VPWR VPWR _2729_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4635_ _1993_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4566_ _0849_ _1955_ _0034_ tree_instances\[4\].u_tree.pipeline_valid\[0\] VGND VGND
+ VPWR VPWR _0162_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_71_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6305_ clknet_leaf_14_clk _0114_ net29 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3517_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1039_ sky130_fd_sc_hd__clkbuf_1
X_4497_ _1902_ _1918_ tree_instances\[8\].u_tree.u_tree_weight_rom.cache_valid VGND
+ VGND VPWR VPWR _0130_ sky130_fd_sc_hd__a21o_1
X_3448_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _0978_ sky130_fd_sc_hd__clkbuf_1
X_6236_ _3117_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__clkbuf_1
X_3379_ _0913_ _0915_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__nor2_1
X_6167_ _3074_ VGND VGND VPWR VPWR _3075_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6801__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5118_ _2305_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__clkbuf_1
X_6098_ tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[2\] _2595_ _0034_ VGND
+ VGND VPWR VPWR _3029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5049_ _1673_ _2221_ VGND VGND VPWR VPWR _2268_ sky130_fd_sc_hd__and2_1
XFILLER_0_94_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4217__B _0799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_75_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5736__A1_N _2708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6542__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4420_ _0977_ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4351_ _1809_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__inv_2
X_4282_ _1743_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__clkbuf_1
X_3302_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[7\] _0846_ VGND VGND
+ VPWR VPWR _0847_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_3_3__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3233_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__clkbuf_1
X_6021_ tree_instances\[3\].u_tree.frame_id_out\[0\] tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0799_ VGND VGND VPWR VPWR _2973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3164_ _0713_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__or2_1
X_6923_ clknet_leaf_73_clk _0636_ net39 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_6854_ clknet_leaf_66_clk _0574_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[2\].u_tree.frame_id_out\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3997_ _1464_ _1475_ _0883_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a21o_1
X_5805_ _2841_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__clkbuf_1
X_6785_ clknet_leaf_7_clk _0519_ net25 VGND VGND VPWR VPWR current_voting_frame\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_259 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5736_ _2708_ tree_instances\[14\].u_tree.frame_id_out\[4\] tree_instances\[14\].u_tree.frame_id_out\[2\]
+ _2714_ VGND VGND VPWR VPWR _2781_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__7000__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5667_ tree_instances\[2\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2712_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4618_ _1983_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_20_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5703__A2 _2583_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5598_ _2598_ tree_instances\[1\].u_tree.frame_id_out\[0\] tree_instances\[1\].u_tree.frame_id_out\[3\]
+ _2606_ _2647_ VGND VGND VPWR VPWR _2648_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_13_540 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4549_ _1947_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6219_ tree_instances\[5\].u_tree.frame_id_out\[3\] tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0903_ VGND VGND VPWR VPWR _3106_ sky130_fd_sc_hd__mux2_1
XANTENNA__5467__A1 _2125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5612__A _2610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_86_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_56_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_97_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkload19 clknet_leaf_9_clk VGND VGND VPWR VPWR clkload19/Y sky130_fd_sc_hd__clkinv_2
XFILLER_0_50_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6723__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_381 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3920_ _1399_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3851_ _1188_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND
+ VPWR VPWR _1336_ sky130_fd_sc_hd__and2b_1
X_3782_ _1262_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6570_ clknet_leaf_61_clk _0339_ net35 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5521_ _2579_ VGND VGND VPWR VPWR _2580_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5452_ _2537_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5697__A1 _2603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6464__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4403_ _1841_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5697__B2 _2659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5383_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[5\] _1247_ VGND VGND
+ VPWR VPWR _2485_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4334_ _1786_ VGND VGND VPWR VPWR _1800_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4747__S _0008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4265_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1733_ sky130_fd_sc_hd__clkbuf_1
X_6004_ tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[0\] _1826_ _0032_ VGND
+ VGND VPWR VPWR _2962_ sky130_fd_sc_hd__mux2_1
X_3216_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0766_ sky130_fd_sc_hd__clkbuf_1
X_4196_ _1661_ VGND VGND VPWR VPWR _1668_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_212 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6906_ clknet_leaf_72_clk _0619_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_25_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6837_ clknet_leaf_79_clk _0557_ net39 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_81_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6768_ clknet_leaf_11_clk _0502_ net25 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.frame_id_in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6699_ clknet_leaf_55_clk _0448_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5719_ _2738_ _2745_ _2755_ _2763_ VGND VGND VPWR VPWR _2764_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5607__A _2578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_92_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5860__A1 _1834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5517__A _2576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4050_ _1504_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3500__A _0733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5603__B2 tree_instances\[1\].u_tree.prediction_out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4952_ _2212_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_1
X_3903_ _1366_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_19_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4883_ _0967_ VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__clkbuf_1
X_6622_ clknet_leaf_58_clk _0381_ net37 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_50_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3834_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1319_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6645__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3765_ _1256_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6553_ clknet_leaf_102_clk _0327_ net32 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_378 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5504_ _2568_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_30_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3696_ _1197_ _1198_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__or2b_1
X_6484_ clknet_leaf_10_clk _0090_ net27 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5435_ _1489_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[6\] _2518_
+ VGND VGND VPWR VPWR _2526_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5366_ _2467_ VGND VGND VPWR VPWR _2468_ sky130_fd_sc_hd__clkbuf_1
X_5297_ _1137_ _2420_ _0016_ tree_instances\[15\].u_tree.pipeline_valid\[0\] VGND
+ VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o2bb2a_1
X_4317_ _1783_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_58_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4248_ _1031_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4179_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1651_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_2_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XPHY_EDGE_ROW_14_Right_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6386__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6315__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5337__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_103_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5530__A0 _2586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_23_Right_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_1_Left_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_32_Right_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6010__A1 _1834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3550_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3481_ _1005_ _1007_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__nor2_1
X_5220_ tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[3\] _2249_ _0020_ VGND
+ VGND VPWR VPWR _2381_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_41_Right_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_47_Left_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5151_ _2324_ VGND VGND VPWR VPWR _2325_ sky130_fd_sc_hd__clkbuf_1
X_5082_ _1547_ _2255_ VGND VGND VPWR VPWR _2285_ sky130_fd_sc_hd__and2_1
X_4102_ _1576_ VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__clkbuf_1
X_4033_ _1509_ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_69_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_56_Left_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_50_Right_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_63_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_35_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5984_ _2950_ VGND VGND VPWR VPWR _2951_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6826__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4935_ _1708_ _2133_ VGND VGND VPWR VPWR _2204_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4866_ _2142_ VGND VGND VPWR VPWR _2147_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6605_ clknet_leaf_36_clk _0369_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3817_ _1009_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4797_ _1698_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[3\] VGND
+ VGND VPWR VPWR _2100_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6536_ clknet_leaf_102_clk _0310_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_3748_ _1241_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6563__SET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6467_ clknet_leaf_28_clk _0255_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_65_Left_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3679_ _1176_ _1181_ _1184_ _0756_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__o31a_1
X_5418_ _1465_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[5\] tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ _1461_ _2514_ VGND VGND VPWR VPWR _2515_ sky130_fd_sc_hd__o221a_1
X_6398_ clknet_leaf_52_clk _0200_ net37 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_370 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5349_ _2449_ _2450_ VGND VGND VPWR VPWR _2451_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_7_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5815__A1 _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_74_Left_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap24 net25 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_12
XFILLER_0_65_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6567__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_50_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_162 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_83_Left_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_571 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6990__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_60_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4720_ _2053_ VGND VGND VPWR VPWR _2054_ sky130_fd_sc_hd__clkbuf_1
X_4651_ tree_instances\[10\].u_tree.read_enable _2008_ VGND VGND VPWR VPWR _2009_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3602_ tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_12_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4582_ _1964_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3533_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6321_ clknet_leaf_84_clk _0129_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[8\].u_tree.pipeline_prediction\[0\]\[0\] sky130_fd_sc_hd__dfrtp_1
X_3464_ tree_instances\[1\].u_tree.ready_for_next tree_instances\[0\].u_tree.ready_for_next
+ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__nand3_1
X_6252_ net13 VGND VGND VPWR VPWR _3125_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6183_ _1888_ _3035_ VGND VGND VPWR VPWR _3087_ sky130_fd_sc_hd__and2_1
X_5203_ _2336_ _2367_ VGND VGND VPWR VPWR _2372_ sky130_fd_sc_hd__and2_1
X_3395_ _0732_ tree_instances\[6\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _0931_ sky130_fd_sc_hd__or2_1
X_5134_ _2315_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5065_ _2276_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__clkbuf_1
X_4016_ _1491_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3284__A1 _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5967_ _0031_ _2934_ VGND VGND VPWR VPWR _2935_ sky130_fd_sc_hd__nor2_1
XANTENNA__6660__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_32_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_4
X_4918_ _1723_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[2\] _2192_
+ VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__mux2_1
X_5898_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_data\[12\] tree_instances\[20\].u_tree.u_tree_weight_rom.gen_tree_20.u_tree_rom.node_data\[12\]
+ _2897_ VGND VGND VPWR VPWR _2898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4849_ _2135_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6519_ clknet_leaf_8_clk _0302_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_99_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_89_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_23_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA__6330__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_91_Left_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5525__A _2582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ tree_instances\[14\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__buf_2
XFILLER_0_28_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6489__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6418__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_62_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6870_ clknet_leaf_78_clk _0589_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_44_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5821_ tree_instances\[0\].u_tree.frame_id_out\[2\] tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0737_ VGND VGND VPWR VPWR _2849_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_17_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5752_ _2583_ _2794_ _2795_ _2796_ tree_instances\[11\].u_tree.prediction_valid VGND
+ VGND VPWR VPWR _2797_ sky130_fd_sc_hd__o221a_1
XANTENNA__5963__B1 _0040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_4
X_4703_ _1590_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND
+ VGND VPWR VPWR _2038_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5683_ _2711_ _2718_ _2635_ _2727_ VGND VGND VPWR VPWR _2728_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_77_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4634_ tree_instances\[10\].u_tree.pipeline_prediction\[0\]\[0\] _1990_ _1992_ VGND
+ VGND VPWR VPWR _1993_ sky130_fd_sc_hd__mux2_1
XANTENNA__4518__A1 _1832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4565_ tree_instances\[4\].u_tree.tree_state\[0\] _0848_ VGND VGND VPWR VPWR _1955_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6304_ clknet_leaf_14_clk _0113_ net30 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3516_ _1035_ _1037_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_4_Right_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4496_ _1917_ VGND VGND VPWR VPWR _1918_ sky130_fd_sc_hd__clkbuf_1
X_3447_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _0977_ sky130_fd_sc_hd__clkbuf_1
X_6235_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[0\] _2456_ _3116_
+ VGND VGND VPWR VPWR _3117_ sky130_fd_sc_hd__mux2_1
X_3378_ _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__clkbuf_1
X_6166_ _3073_ VGND VGND VPWR VPWR _3074_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5117_ tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[0\] _2122_ _0018_ VGND
+ VGND VPWR VPWR _2305_ sky130_fd_sc_hd__mux2_1
X_6097_ _3028_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__clkbuf_1
X_5048_ _2267_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6841__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6999_ clknet_leaf_51_clk _0065_ net35 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_82_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6929__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4395__S _0040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6582__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6511__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_14_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_207 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4350_ _1803_ tree_instances\[16\].u_tree.pipeline_valid\[0\] tree_instances\[16\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__or3b_2
XFILLER_0_111_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3301_ _0845_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__clkbuf_1
X_4281_ _1748_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__clkbuf_1
X_3232_ _0780_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_3_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_4
X_6020_ _2969_ _2970_ _2972_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__o21ai_1
X_3163_ _0714_ _0718_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__or2_1
XANTENNA__5702__B _2588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6922_ clknet_leaf_74_clk _0635_ net39 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6853_ clknet_leaf_40_clk _0573_ net30 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4739__A1 _1827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5804_ _2839_ _2840_ VGND VGND VPWR VPWR _2841_ sky130_fd_sc_hd__and2_1
XANTENNA__6025__S _0799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3996_ _1468_ _1474_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__nor2_1
X_6784_ clknet_leaf_7_clk _0518_ net25 VGND VGND VPWR VPWR current_voting_frame\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5735_ _2773_ _2774_ _2779_ VGND VGND VPWR VPWR _2780_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5666_ _2708_ tree_instances\[2\].u_tree.frame_id_out\[4\] _2710_ VGND VGND VPWR
+ VPWR _2711_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_44_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4617_ _1788_ _1937_ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_20_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5597_ _2578_ tree_instances\[1\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2647_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4548_ _1742_ _1945_ VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4479_ tree_instances\[8\].u_tree.read_enable VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__clkbuf_1
X_6218_ _3105_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__clkbuf_1
X_6149_ _2176_ _2179_ _2183_ _2184_ VGND VGND VPWR VPWR _3060_ sky130_fd_sc_hd__or4_1
XTAP_TAPCELL_ROW_86_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_79_Right_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_56_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_97_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_88_Right_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5803__A _2586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6763__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Right_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_98_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_106_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3850_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1335_ sky130_fd_sc_hd__inv_2
X_3781_ _1270_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5520_ _2578_ VGND VGND VPWR VPWR _2579_ sky130_fd_sc_hd__clkbuf_4
X_5451_ _1494_ _2534_ VGND VGND VPWR VPWR _2537_ sky130_fd_sc_hd__and2_1
XANTENNA__5146__B2 tree_instances\[16\].u_tree.ready_for_next VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_4402_ tree_instances\[7\].u_tree.frame_id_out\[0\] tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0970_ VGND VGND VPWR VPWR _1841_ sky130_fd_sc_hd__mux2_1
X_5382_ _2483_ VGND VGND VPWR VPWR _2484_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5720__A1_N _2708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4333_ _1795_ VGND VGND VPWR VPWR _1799_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5713__A _2622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4264_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1732_ sky130_fd_sc_hd__clkbuf_1
X_3215_ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__clkbuf_1
X_6003_ _2961_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4195_ _1660_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__clkbuf_1
X_6905_ clknet_leaf_72_clk _0618_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_10_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_53_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6836_ clknet_leaf_84_clk _0556_ net39 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_81_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6767_ clknet_leaf_11_clk _0501_ net25 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.frame_id_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3979_ _1458_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
X_5718_ _2713_ tree_instances\[18\].u_tree.frame_id_out\[1\] _2756_ _2762_ tree_instances\[18\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2763_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_33_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6698_ clknet_leaf_55_clk _0447_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5649_ state\[0\] _2447_ attack_votes\[1\] VGND VGND VPWR VPWR _2698_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5623__A _2585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_92_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_5_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6944__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5533__A _2588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5300__A1 _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4951_ _1827_ tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[0\] _1824_ VGND
+ VGND VPWR VPWR _2212_ sky130_fd_sc_hd__mux2_1
X_3902_ _0913_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4882_ _2158_ VGND VGND VPWR VPWR _2163_ sky130_fd_sc_hd__clkbuf_1
X_6621_ clknet_leaf_34_clk _0380_ VGND VGND VPWR VPWR tree_instances\[16\].u_tree.u_tree_weight_rom.cached_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_50_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3833_ _1191_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6552_ clknet_leaf_45_clk _0326_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3764_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_485 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5119__A1 _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5503_ _2478_ _2484_ _2493_ VGND VGND VPWR VPWR _2568_ sky130_fd_sc_hd__and3_1
X_6483_ clknet_leaf_9_clk _0271_ net27 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XTAP_TAPCELL_ROW_30_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3695_ _0731_ tree_instances\[20\].u_tree.pipeline_valid\[0\] tree_instances\[20\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__o21ai_1
X_5434_ _2525_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6685__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_538 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6614__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5365_ _2448_ VGND VGND VPWR VPWR _2467_ sky130_fd_sc_hd__clkbuf_1
X_5296_ tree_instances\[15\].u_tree.pipeline_valid\[0\] tree_instances\[15\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _2420_ sky130_fd_sc_hd__nand2_1
X_4316_ _1035_ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_58_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4247_ _1715_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__clkbuf_1
X_4178_ _1649_ VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__buf_1
XFILLER_0_97_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_2_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_66_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6424__D _0032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6819_ clknet_leaf_52_clk _0540_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_94_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_94_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6355__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_103_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_352 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_max_cap26_A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3480_ _1006_ tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND
+ VPWR VPWR _1007_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_102_Left_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _0786_ VGND VGND VPWR VPWR _2324_ sky130_fd_sc_hd__clkbuf_1
X_5081_ _2284_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__clkbuf_1
X_4101_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1576_ sky130_fd_sc_hd__clkbuf_1
X_4032_ _1508_ VGND VGND VPWR VPWR _1509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_69_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5983_ _2949_ VGND VGND VPWR VPWR _2950_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_111_Left_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_63_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4934_ _2203_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_35_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4865_ _0813_ VGND VGND VPWR VPWR _2146_ sky130_fd_sc_hd__clkbuf_1
X_3816_ _1297_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__clkbuf_1
X_6604_ clknet_leaf_39_clk _0368_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4796_ _2094_ _2095_ _2096_ _2097_ _2098_ VGND VGND VPWR VPWR _2099_ sky130_fd_sc_hd__a221o_1
XANTENNA__6866__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3747_ _1240_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND
+ VPWR VPWR _1241_ sky130_fd_sc_hd__nor2_1
X_6535_ clknet_leaf_1_clk _0309_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_6466_ clknet_leaf_27_clk _0254_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3678_ _1182_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5417_ _0868_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[3\] VGND
+ VGND VPWR VPWR _2514_ sky130_fd_sc_hd__xnor2_1
X_6397_ clknet_leaf_52_clk _0199_ net35 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5348_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _2450_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_7_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5279_ tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[3\] _2249_ _0022_ VGND
+ VGND VPWR VPWR _2411_ sky130_fd_sc_hd__mux2_1
Xmax_cap25 net27 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__buf_12
XFILLER_0_97_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5579__A1 _2575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5551__A1_N _2598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_366 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4398__S _0040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_12 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_32_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4650_ _1998_ _2001_ _2005_ _2007_ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__or4_1
X_3601_ tree_instances\[0\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5742__A1 _2709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6320_ clknet_leaf_56_clk _0128_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_12_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4581_ _1764_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[6\] _1956_
+ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3532_ _1052_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3463_ tree_instances\[3\].u_tree.ready_for_next tree_instances\[2\].u_tree.ready_for_next
+ tree_instances\[5\].u_tree.ready_for_next tree_instances\[4\].u_tree.ready_for_next
+ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6251_ _2998_ _3010_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__nor2_1
X_6182_ _3086_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__clkbuf_1
X_5202_ _2371_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__clkbuf_1
X_3394_ _0912_ _0918_ _0924_ _0930_ tree_instances\[16\].u_tree.tree_state\[1\] VGND
+ VGND VPWR VPWR _0060_ sky130_fd_sc_hd__a41o_1
X_5133_ tree_instances\[16\].u_tree.frame_id_out\[0\] tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _1023_ VGND VGND VPWR VPWR _2315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5064_ tree_instances\[15\].u_tree.frame_id_out\[0\] tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _1137_ VGND VGND VPWR VPWR _2276_ sky130_fd_sc_hd__mux2_1
X_4015_ _1485_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_406 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_48_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5966_ tree_instances\[3\].u_tree.tree_state\[0\] _0850_ tree_instances\[3\].u_tree.tree_state\[1\]
+ _0800_ VGND VGND VPWR VPWR _2934_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_74_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4917_ _2194_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__clkbuf_1
X_5897_ _2896_ VGND VGND VPWR VPWR _2897_ sky130_fd_sc_hd__clkbuf_1
X_4848_ tree_instances\[12\].u_tree.frame_id_out\[1\] tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0829_ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4779_ tree_instances\[11\].u_tree.tree_state\[3\] _0952_ _1816_ tree_instances\[11\].u_tree.ready_for_next
+ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__a22o_1
XANTENNA__5733__A1 _2627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5733__B2 _2619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6518_ clknet_leaf_8_clk _0301_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6449_ clknet_leaf_97_clk _0242_ net32 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5631__A _2582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_89_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6788__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5724__B2 _2598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5806__A _2589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6370__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_509 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_111_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5541__A _1832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_109_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5820_ _2848_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_17_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5751_ _2589_ tree_instances\[11\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2796_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__6458__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4702_ _1591_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND
+ VGND VPWR VPWR _2037_ sky130_fd_sc_hd__nand2_1
X_5682_ _2583_ _2719_ tree_instances\[4\].u_tree.prediction_valid _2720_ _2726_ VGND
+ VGND VPWR VPWR _2727_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_71_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4633_ tree_instances\[10\].u_tree.tree_state\[0\] tree_instances\[10\].u_tree.tree_state\[1\]
+ tree_instances\[10\].u_tree.tree_state\[2\] _1991_ _1170_ VGND VGND VPWR VPWR _1992_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_25_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_77_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4564_ _1954_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6303_ clknet_leaf_19_clk _0112_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3515_ _1036_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4495_ _1908_ _1912_ _1914_ _1916_ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__or4_2
X_6234_ net15 VGND VGND VPWR VPWR _3116_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_110_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3446_ _0975_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3377_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _0914_ sky130_fd_sc_hd__clkbuf_1
X_6165_ _0717_ VGND VGND VPWR VPWR _3073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6096_ tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[1\] _1829_ _0034_ VGND
+ VGND VPWR VPWR _3028_ sky130_fd_sc_hd__mux2_1
X_5116_ _2304_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__clkbuf_1
X_5047_ _1669_ _2222_ VGND VGND VPWR VPWR _2267_ sky130_fd_sc_hd__and2_1
XFILLER_0_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6998_ clknet_leaf_38_clk _0104_ net29 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6881__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5949_ _1431_ _2553_ VGND VGND VPWR VPWR _2925_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_14_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6551__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3300_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _0845_ sky130_fd_sc_hd__buf_1
X_4280_ _1740_ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__clkbuf_1
X_3231_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0780_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3162_ _0715_ _0716_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_72_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6639__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6921_ clknet_leaf_73_clk _0634_ net39 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6852_ clknet_leaf_66_clk _0572_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[2\].u_tree.frame_id_out\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5803_ _2586_ _2837_ VGND VGND VPWR VPWR _2840_ sky130_fd_sc_hd__or2_1
X_3995_ _1470_ _1473_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6783_ clknet_leaf_19_clk _0517_ net25 VGND VGND VPWR VPWR current_voting_frame\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5734_ _2709_ tree_instances\[19\].u_tree.frame_id_out\[3\] _2775_ _2778_ VGND VGND
+ VPWR VPWR _2779_ sky130_fd_sc_hd__o211a_1
XFILLER_0_72_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5665_ _2709_ tree_instances\[2\].u_tree.frame_id_out\[3\] tree_instances\[2\].u_tree.frame_id_out\[4\]
+ _2708_ VGND VGND VPWR VPWR _2710_ sky130_fd_sc_hd__o22a_1
XFILLER_0_32_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4350__A _1803_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4616_ _1982_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_111_Right_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5596_ _2583_ tree_instances\[1\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2646_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4547_ _1946_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4478_ _1900_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
X_3429_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _0962_ sky130_fd_sc_hd__inv_2
X_6217_ tree_instances\[5\].u_tree.frame_id_out\[2\] tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0903_ VGND VGND VPWR VPWR _3105_ sky130_fd_sc_hd__mux2_1
X_6148_ _1686_ _2170_ _3057_ _3058_ _2169_ VGND VGND VPWR VPWR _3059_ sky130_fd_sc_hd__a221o_1
X_6079_ _3018_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_86_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_56_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_28_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6309__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5927__A1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_97_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_61_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_76_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6732__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3780_ _1265_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_14_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5450_ _2536_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4401_ _1839_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_1_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_29_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5381_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[7\] _2473_ VGND VGND
+ VPWR VPWR _2483_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4332_ _1798_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4263_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1731_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3214_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _0764_ sky130_fd_sc_hd__clkbuf_1
X_6002_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[7\] _1425_ _2959_
+ VGND VGND VPWR VPWR _2961_ sky130_fd_sc_hd__mux2_1
X_4194_ _1664_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6473__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6904_ clknet_leaf_72_clk _0617_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_77_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_53_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_25_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6402__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6835_ clknet_leaf_74_clk _0555_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.cached_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3978_ tree_instances\[16\].u_tree.prediction_valid _1023_ VGND VGND VPWR VPWR _1458_
+ sky130_fd_sc_hd__and2b_1
X_6766_ clknet_leaf_11_clk _0500_ net24 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.frame_id_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5717_ _2619_ tree_instances\[18\].u_tree.frame_id_out\[2\] _2757_ _2586_ _2761_
+ VGND VGND VPWR VPWR _2762_ sky130_fd_sc_hd__o221a_1
X_6697_ clknet_leaf_54_clk _0446_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5648_ _2693_ _2614_ VGND VGND VPWR VPWR _2697_ sky130_fd_sc_hd__or2b_1
X_5579_ _2575_ tree_instances\[3\].u_tree.frame_id_out\[0\] tree_instances\[3\].u_tree.frame_id_out\[1\]
+ _2602_ VGND VGND VPWR VPWR _2629_ sky130_fd_sc_hd__o22a_1
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_92_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_5_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_570 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6984__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6913__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4950_ _2211_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__clkbuf_1
X_3901_ _1377_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4881_ _2155_ VGND VGND VPWR VPWR _2162_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6620_ clknet_leaf_20_clk _0086_ net25 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3832_ _1195_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_50_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6551_ clknet_leaf_44_clk _0325_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5502_ _2566_ VGND VGND VPWR VPWR _2567_ sky130_fd_sc_hd__clkbuf_1
X_3763_ _0745_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5772__C1 _2613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_114 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6482_ clknet_leaf_98_clk _0270_ net27 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.prediction_out
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3694_ tree_instances\[20\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__buf_2
XFILLER_0_42_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5433_ _1480_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[5\] _2518_
+ VGND VGND VPWR VPWR _2525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5364_ _2458_ VGND VGND VPWR VPWR _2466_ sky130_fd_sc_hd__clkbuf_1
X_4315_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1782_ sky130_fd_sc_hd__inv_2
X_5295_ _0753_ _1884_ _1801_ tree_instances\[18\].u_tree.ready_for_next VGND VGND
+ VPWR VPWR _0429_ sky130_fd_sc_hd__a22o_1
X_4246_ _1714_ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6654__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_58_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4177_ _1648_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5055__A1 _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6818_ clknet_leaf_52_clk _0539_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4566__B1 _0034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6749_ clknet_leaf_98_clk _0005_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5337__C _0996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_94_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6395__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6324__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_139 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5544__A _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5080_ _1544_ _2255_ VGND VGND VPWR VPWR _2284_ sky130_fd_sc_hd__and2_1
X_4100_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1575_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4031_ _1507_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_69_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5982_ _2948_ VGND VGND VPWR VPWR _2949_ sky130_fd_sc_hd__buf_1
XFILLER_0_63_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4933_ _1673_ _1683_ _1685_ VGND VGND VPWR VPWR _2203_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_35_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4864_ _2144_ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__clkbuf_1
X_6603_ clknet_leaf_38_clk _0367_ net30 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3815_ _1303_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4795_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[6\] tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__xor2_1
XFILLER_0_104_108 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3746_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1240_ sky130_fd_sc_hd__buf_1
X_6534_ clknet_leaf_0_clk _0308_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_6465_ clknet_leaf_28_clk _0253_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5416_ _1471_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[2\] tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ _1465_ VGND VGND VPWR VPWR _2513_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3677_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[3\] _0766_ VGND VGND
+ VPWR VPWR _1183_ sky130_fd_sc_hd__nor2_1
X_6396_ clknet_leaf_52_clk _0198_ net35 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5347_ _1240_ VGND VGND VPWR VPWR _2449_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_7_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5278_ _2410_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__clkbuf_1
X_4229_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1698_ sky130_fd_sc_hd__inv_2
Xmax_cap15 net16 VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
Xmax_cap26 net32 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__buf_12
XFILLER_0_65_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6576__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6505__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5019__A1 _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_24 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_610 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_60_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3600_ _1058_ _1067_ _1051_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a21boi_1
X_4580_ _1963_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3531_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1052_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_12_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_110_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3462_ _0971_ _0988_ _0991_ tree_instances\[6\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0080_ sky130_fd_sc_hd__a31o_1
X_6250_ _3124_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3393_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__clkbuf_1
X_6181_ _3076_ _3035_ VGND VGND VPWR VPWR _3086_ sky130_fd_sc_hd__and2_1
X_5201_ _2332_ _2367_ VGND VGND VPWR VPWR _2371_ sky130_fd_sc_hd__and2_1
X_5132_ _2311_ _2312_ _2314_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__o21ai_1
X_5063_ _0016_ VGND VGND VPWR VPWR _2275_ sky130_fd_sc_hd__inv_2
X_4014_ _1488_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_48_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5965_ tree_instances\[3\].u_tree.tree_state\[1\] tree_instances\[3\].u_tree.current_node_data\[107\]
+ tree_instances\[3\].u_tree.node_data\[107\] _2932_ VGND VGND VPWR VPWR _2933_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4916_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[1\] _1713_ tree_instances\[12\].u_tree.read_enable
+ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__mux2_1
X_5896_ _2895_ VGND VGND VPWR VPWR _2896_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4847_ _2134_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4778_ _2084_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkbuf_1
X_3729_ tree_instances\[1\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__buf_2
X_6517_ clknet_leaf_8_clk _0300_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6448_ clknet_leaf_100_clk _0241_ net32 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6379_ clknet_leaf_81_clk _0186_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_277 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6757__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_100_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_45_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5750_ _2588_ tree_instances\[11\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2795_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_84_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5681_ _2627_ _2721_ _2722_ _2723_ _2725_ VGND VGND VPWR VPWR _2726_ sky130_fd_sc_hd__o221a_1
XFILLER_0_60_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4701_ _0829_ _0830_ _0010_ tree_instances\[12\].u_tree.pipeline_valid\[0\] VGND
+ VGND VPWR VPWR _0216_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4632_ tree_instances\[10\].u_tree.tree_state\[0\] _1135_ VGND VGND VPWR VPWR _1991_
+ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_77_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4563_ _1724_ _1701_ _1706_ _1722_ VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6302_ clknet_leaf_13_clk _0111_ net29 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_4494_ _1791_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[1\] tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ _1775_ _1915_ VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__a221o_1
X_3514_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1036_ sky130_fd_sc_hd__buf_1
X_3445_ _0972_ _0974_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__or2_1
X_6233_ _3110_ tree_instances\[16\].u_tree.node_data\[12\] _3115_ VGND VGND VPWR VPWR
+ _0672_ sky130_fd_sc_hd__a21o_1
XANTENNA__5732__A _2579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3376_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _0913_ sky130_fd_sc_hd__buf_1
X_6164_ tree_instances\[20\].u_tree.u_tree_weight_rom.gen_tree_20.u_tree_rom.node_data\[12\]
+ _3068_ _3071_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_data\[12\] _3072_
+ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__a221o_1
X_6095_ _3027_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__clkbuf_1
X_5115_ _1444_ _2296_ VGND VGND VPWR VPWR _2304_ sky130_fd_sc_hd__and2_1
XANTENNA__4348__A _1803_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5046_ _2266_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6997_ clknet_leaf_31_clk _0703_ net29 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
X_5948_ _2924_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5879_ _2880_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6850__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_261 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_14_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6938__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6591__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5536__B _2441_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6520__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3230_ _0778_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__clkbuf_1
X_3161_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _0717_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6920_ clknet_leaf_73_clk _0633_ net39 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_21 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4615__B _1937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6851_ clknet_leaf_74_clk _0571_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.current_node_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_5802_ _2586_ _2837_ VGND VGND VPWR VPWR _2839_ sky130_fd_sc_hd__nand2_1
X_3994_ _1471_ _1472_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_83_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6782_ clknet_leaf_7_clk _0516_ net24 VGND VGND VPWR VPWR current_voting_frame\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5733_ _2627_ _2776_ tree_instances\[19\].u_tree.frame_id_out\[2\] _2619_ _2777_
+ VGND VGND VPWR VPWR _2778_ sky130_fd_sc_hd__o221a_1
XANTENNA__6608__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5664_ _2606_ VGND VGND VPWR VPWR _2709_ sky130_fd_sc_hd__buf_2
X_4615_ _1797_ _1937_ VGND VGND VPWR VPWR _1982_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5595_ _2638_ _2641_ _2644_ VGND VGND VPWR VPWR _2645_ sky130_fd_sc_hd__and3b_1
XFILLER_0_102_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4546_ _1750_ _1945_ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4477_ tree_instances\[8\].u_tree.pipeline_prediction\[0\]\[0\] _1896_ _1899_ VGND
+ VGND VPWR VPWR _1900_ sky130_fd_sc_hd__mux2_1
X_3428_ _0957_ _0960_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__nor2_1
X_6216_ _3104_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__clkbuf_1
X_3359_ _0896_ _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__nand2_1
X_6147_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[6\] tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ VGND VGND VPWR VPWR _3058_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_318 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6078_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[2\] _1350_ _2989_
+ VGND VGND VPWR VPWR _3018_ sky130_fd_sc_hd__mux2_1
X_5029_ tree_instances\[14\].u_tree.frame_id_out\[2\] tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0735_ VGND VGND VPWR VPWR _2258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6349__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_97_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_88_Left_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6772__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6701__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4400_ tree_instances\[7\].u_tree.tree_state\[2\] tree_instances\[7\].u_tree.tree_state\[1\]
+ _1812_ VGND VGND VPWR VPWR _1839_ sky130_fd_sc_hd__or3_1
XFILLER_0_50_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5380_ _2479_ VGND VGND VPWR VPWR _2482_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4331_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[7\] _1796_ _1792_ VGND
+ VGND VPWR VPWR _1798_ sky130_fd_sc_hd__and3_1
X_4262_ _1729_ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5854__A1 _1826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3213_ _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__clkbuf_1
X_6001_ _2960_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__clkbuf_1
X_4193_ _1651_ _0956_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_77_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6903_ clknet_leaf_73_clk _0616_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6834_ clknet_leaf_40_clk _0098_ net30 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
X_6765_ clknet_leaf_26_clk _0499_ net24 VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__dfrtp_1
X_3977_ _1450_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__clkbuf_1
X_5716_ _2606_ tree_instances\[18\].u_tree.frame_id_out\[3\] _2758_ _2759_ _2760_
+ VGND VGND VPWR VPWR _2761_ sky130_fd_sc_hd__o221a_1
XANTENNA__6442__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4593__A1 _1832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6696_ clknet_leaf_54_clk _0445_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_487 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5647_ _2690_ _2693_ _2695_ attack_votes\[1\] VGND VGND VPWR VPWR _2696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5578_ tree_instances\[3\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2628_ sky130_fd_sc_hd__inv_2
XANTENNA__5542__B1 _1835_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4529_ _1936_ VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6098__A1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_5_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_80_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6261__A1 _1834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6953__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3900_ _1381_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_4
X_4880_ _2148_ VGND VGND VPWR VPWR _2161_ sky130_fd_sc_hd__clkbuf_1
X_3831_ _1316_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
X_3762_ _1253_ _0742_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_80_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6550_ clknet_leaf_42_clk _0324_ net36 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5501_ _0714_ VGND VGND VPWR VPWR _2566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6481_ clknet_leaf_92_clk _0269_ net27 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_30_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3693_ _0809_ _0828_ _0802_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__a21boi_1
X_5432_ _2524_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__clkbuf_1
X_5363_ _2459_ VGND VGND VPWR VPWR _2465_ sky130_fd_sc_hd__buf_1
XFILLER_0_77_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4314_ _1780_ VGND VGND VPWR VPWR _1781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5294_ _2419_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__clkbuf_1
X_4245_ _1697_ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_58_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4176_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1648_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4356__A _1803_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6694__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_2_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_2_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6623__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_62_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_60_clk_A clknet_3_7__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6004__A1 _1826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6817_ clknet_leaf_53_clk _0538_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output8_A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6748_ clknet_leaf_92_clk _0047_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_33_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6679_ clknet_leaf_56_clk _0429_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_60_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_103_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5754__B1 _2798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5544__B _1834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5809__A1 _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4030_ _0898_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_10_Right_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_16_Left_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5981_ tree_instances\[3\].u_tree.read_enable _2947_ VGND VGND VPWR VPWR _2948_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_44_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_4
X_4932_ _2202_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_35_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_63_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6602_ clknet_leaf_39_clk _0366_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4623__B _1937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_25_Left_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4863_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _2144_ sky130_fd_sc_hd__clkbuf_1
X_3814_ _1291_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4342__C net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4794_ _0837_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[1\] VGND
+ VGND VPWR VPWR _2097_ sky130_fd_sc_hd__or2_1
X_3745_ _0789_ _1237_ _1239_ _0776_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__o31a_1
XFILLER_0_15_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6533_ clknet_leaf_102_clk _0307_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_6464_ clknet_leaf_27_clk _0252_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5415_ _1461_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[6\] tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ _1459_ VGND VGND VPWR VPWR _2512_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3676_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[1\] tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[0\]
+ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6395_ clknet_leaf_52_clk _0197_ net37 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_7_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5346_ _0938_ VGND VGND VPWR VPWR _2448_ sky130_fd_sc_hd__clkbuf_1
X_5277_ tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[2\] _2125_ _0022_ VGND
+ VGND VPWR VPWR _2410_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_34_Left_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4228_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1697_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6804__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4159_ _1630_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_106_Right_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xmax_cap16 net41 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
Xmax_cap27 net32 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__buf_12
XFILLER_0_78_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_35_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_93_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_43_Left_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_52_Left_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6545__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_load_slew38_A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_61_Left_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_26_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_84_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_32_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_60_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_154 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_368 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3530_ tree_instances\[15\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_12_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3461_ _0989_ _0990_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__nor2_1
XPHY_EDGE_ROW_70_Left_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3392_ _0928_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__clkbuf_1
X_5200_ _2370_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__clkbuf_1
X_6180_ tree_instances\[5\].u_tree.u_tree_weight_rom.cache_valid _3011_ _3010_ VGND
+ VGND VPWR VPWR _0649_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_460 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5131_ _2313_ VGND VGND VPWR VPWR _2314_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_20_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5062_ _2274_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__clkbuf_1
X_4013_ _0872_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_3_6__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6207__A1 tree_instances\[0\].u_tree.frame_id_in\[4\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__4337__C net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_48_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_482 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_17_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5964_ _0850_ VGND VGND VPWR VPWR _2932_ sky130_fd_sc_hd__clkbuf_1
X_4915_ _2193_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_1
X_5895_ _2894_ tree_instances\[20\].u_tree.read_enable VGND VGND VPWR VPWR _2895_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4846_ tree_instances\[12\].u_tree.frame_id_out\[0\] tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0829_ VGND VGND VPWR VPWR _2134_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4777_ _1604_ _2029_ VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__and2_1
X_6516_ clknet_leaf_7_clk _0299_ net25 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3728_ _0731_ tree_instances\[1\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _1226_ sky130_fd_sc_hd__or2_1
XANTENNA__7003__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3659_ _1167_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__clkbuf_1
X_6447_ clknet_leaf_96_clk _0240_ net32 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6378_ clknet_leaf_80_clk _0185_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_167 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5329_ _2437_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6797__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_111_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6726__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3623__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_109_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_66_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _2576_ tree_instances\[4\].u_tree.frame_id_out\[0\] tree_instances\[4\].u_tree.frame_id_out\[2\]
+ _2714_ _2724_ VGND VGND VPWR VPWR _2725_ sky130_fd_sc_hd__o221a_1
X_4700_ _1136_ _1991_ _1819_ tree_instances\[10\].u_tree.ready_for_next VGND VGND
+ VPWR VPWR _0215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4631_ tree_instances\[10\].u_tree.tree_state\[1\] tree_instances\[10\].u_tree.current_node_data\[12\]
+ tree_instances\[10\].u_tree.node_data\[12\] _1171_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4562_ _1197_ _1198_ _0028_ tree_instances\[20\].u_tree.pipeline_valid\[0\] VGND
+ VGND VPWR VPWR _0160_ sky130_fd_sc_hd__o2bb2a_1
X_6301_ clknet_leaf_40_clk _0110_ net30 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4493_ _1775_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[5\] tree_instances\[8\].u_tree.u_tree_weight_rom.cache_valid
+ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__o21ai_1
X_3513_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6232_ tree_instances\[16\].u_tree.u_tree_weight_rom.gen_tree_16.u_tree_rom.node_data\[12\]
+ _3111_ _3114_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_data\[12\] VGND
+ VGND VPWR VPWR _3115_ sky130_fd_sc_hd__a22o_1
X_3444_ _0973_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_6_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA__6467__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3375_ tree_instances\[16\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__clkbuf_1
X_6163_ _2502_ tree_instances\[20\].u_tree.node_data\[12\] VGND VGND VPWR VPWR _3072_
+ sky130_fd_sc_hd__and2b_1
X_6094_ tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[0\] _1826_ _0034_ VGND
+ VGND VPWR VPWR _3027_ sky130_fd_sc_hd__mux2_1
X_5114_ _2303_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_108_Left_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5045_ _1676_ _2222_ VGND VGND VPWR VPWR _2266_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_88_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_202 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4364__A _1112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6996_ clknet_leaf_83_clk _0702_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5947_ _1422_ _2553_ VGND VGND VPWR VPWR _2924_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5878_ tree_instances\[1\].u_tree.prediction_out tree_instances\[1\].u_tree.pipeline_prediction\[0\]\[0\]
+ tree_instances\[1\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4829_ tree_instances\[12\].u_tree.pipeline_frame_id\[0\]\[0\] _2122_ _0010_ VGND
+ VGND VPWR VPWR _2123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6529__SET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_42_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6978__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_22_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6560__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3160_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _0716_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_72_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6850_ clknet_leaf_67_clk _0570_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5801_ _2837_ _2838_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__nor2_1
X_6781_ clknet_leaf_7_clk _0515_ net25 VGND VGND VPWR VPWR current_voting_frame\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_9_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_8_Right_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3993_ _0867_ _0870_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__nand2_1
X_5732_ _2579_ tree_instances\[19\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2777_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_77 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5663_ _2631_ VGND VGND VPWR VPWR _2708_ sky130_fd_sc_hd__buf_2
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4614_ _1981_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
X_5594_ _2599_ tree_instances\[13\].u_tree.frame_id_out\[2\] _2642_ _2643_ tree_instances\[13\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2644_ sky130_fd_sc_hd__o221a_1
XANTENNA__6648__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4545_ _1944_ VGND VGND VPWR VPWR _1945_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4476_ _0041_ _1898_ VGND VGND VPWR VPWR _1899_ sky130_fd_sc_hd__nor2_1
X_3427_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_39_Right_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6215_ tree_instances\[5\].u_tree.frame_id_out\[1\] tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0903_ VGND VGND VPWR VPWR _3104_ sky130_fd_sc_hd__mux2_1
X_3358_ _0897_ _0898_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__nor2_1
X_6146_ _1661_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[6\] VGND
+ VGND VPWR VPWR _3057_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3289_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _0834_ sky130_fd_sc_hd__clkbuf_1
X_6077_ _3017_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5648__B_N _2614_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5028_ _2257_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6979_ clknet_leaf_38_clk _0685_ net29 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_48_Right_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3438__A _0733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6389__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6790__SET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_57_Right_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_106_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_66_Right_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_55_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5547__B _1020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6741__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_75_Right_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5551__B2 _2600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4330_ _1771_ VGND VGND VPWR VPWR _1797_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4261_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1729_ sky130_fd_sc_hd__clkbuf_1
X_3212_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[1\] tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[0\]
+ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__or2_1
X_6000_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[6\] _1428_ _2959_
+ VGND VGND VPWR VPWR _2960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4192_ _1659_ VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_84_Right_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6902_ clknet_leaf_74_clk _0615_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_6833_ clknet_leaf_46_clk _0554_ net36 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_77_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6764_ clknet_leaf_26_clk _0498_ net24 VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__dfrtp_1
X_3976_ _1449_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6695_ clknet_leaf_57_clk _0444_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6829__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5715_ _2588_ tree_instances\[18\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2760_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__5790__A1 _2820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5646_ _2694_ net11 _2636_ VGND VGND VPWR VPWR _2695_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_93_Right_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6482__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5577_ _2622_ VGND VGND VPWR VPWR _2627_ sky130_fd_sc_hd__buf_4
XANTENNA__5542__A1 _1832_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6411__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4528_ tree_instances\[8\].u_tree.tree_state\[2\] tree_instances\[8\].u_tree.tree_state\[1\]
+ _1813_ VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__or3_1
X_4459_ _0970_ _1883_ _1812_ tree_instances\[7\].u_tree.ready_for_next VGND VGND VPWR
+ VPWR _0127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6129_ _1352_ _2972_ VGND VGND VPWR VPWR _3046_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_24_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_101_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_594 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6993__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3830_ tree_instances\[12\].u_tree.prediction_valid _0829_ VGND VGND VPWR VPWR _1316_
+ sky130_fd_sc_hd__and2b_1
X_3761_ _0746_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_80_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6922__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5500_ _2564_ VGND VGND VPWR VPWR _2565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_338 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3692_ _1186_ _1194_ _1196_ _0850_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__o31a_1
XTAP_TAPCELL_ROW_30_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6480_ clknet_leaf_9_clk _0268_ net27 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5431_ _1495_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[4\] _2519_
+ VGND VGND VPWR VPWR _2524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5362_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _2464_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4313_ _1774_ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6999__SET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_87 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5293_ tree_instances\[18\].u_tree.frame_id_out\[4\] tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[18\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2419_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_91_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4244_ _1703_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__clkbuf_1
X_4175_ _1646_ VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_2_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_66_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_38_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6816_ clknet_leaf_55_clk _0537_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4372__A _1112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6747_ clknet_leaf_82_clk _0490_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.gen_tree_5.u_tree_rom.node_data\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5763__B2 _2606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3959_ _1438_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__clkbuf_1
X_6678_ clknet_leaf_57_clk _0428_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_302 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_94_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5629_ _2673_ _2675_ _2678_ VGND VGND VPWR VPWR _2679_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6333__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_447 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_480 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_69_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6343__SET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5980_ _2937_ _2938_ _2943_ _2946_ VGND VGND VPWR VPWR _2947_ sky130_fd_sc_hd__or4b_1
XFILLER_0_86_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4931_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_data\[12\] tree_instances\[12\].u_tree.u_tree_weight_rom.gen_tree_12.u_tree_rom.node_data\[12\]
+ _2201_ VGND VGND VPWR VPWR _2202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_63_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4862_ _0821_ VGND VGND VPWR VPWR _2143_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_35_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6601_ clknet_leaf_37_clk _0365_ net30 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3813_ _1301_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4793_ _0838_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[1\] VGND
+ VGND VPWR VPWR _2096_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6532_ clknet_leaf_31_clk _0080_ net33 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3744_ _1238_ _0777_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6463_ clknet_leaf_27_clk _0251_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3675_ _1177_ _1180_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5414_ _1482_ _2504_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ _1460_ VGND VGND VPWR VPWR _2511_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_70_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6394_ clknet_leaf_52_clk _0196_ net35 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5751__A _2589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5345_ _2447_ _2445_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_7_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5276_ _2409_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__clkbuf_1
X_4227_ _1695_ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__clkbuf_1
X_4158_ _1626_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__clkbuf_1
Xmax_cap17 _0883_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__buf_1
XFILLER_0_97_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4089_ _1563_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap39 tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_12
XANTENNA__6844__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5736__B2 _2714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6416__SET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6514__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_max_cap24_A net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_12_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_40_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3460_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[7\] tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[6\]
+ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3391_ _0925_ _0927_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__nor2_1
X_5130_ tree_instances\[16\].u_tree.tree_state\[1\] tree_instances\[16\].u_tree.tree_state\[2\]
+ _1809_ VGND VGND VPWR VPWR _2313_ sky130_fd_sc_hd__or3_1
XFILLER_0_58_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5061_ tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[4\] _2251_ _0016_ VGND
+ VGND VPWR VPWR _2274_ sky130_fd_sc_hd__mux2_1
X_4012_ _0876_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5963_ _0970_ _2931_ _0040_ tree_instances\[7\].u_tree.pipeline_valid\[0\] VGND VGND
+ VPWR VPWR _0586_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_48_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4914_ _1708_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[0\] _2192_
+ VGND VGND VPWR VPWR _2193_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_314 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_87_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5894_ _2884_ _2886_ _2893_ VGND VGND VPWR VPWR _2894_ sky130_fd_sc_hd__and3b_1
XANTENNA_clkbuf_leaf_89_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_155 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5718__A1 _2713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4845_ _2130_ _2131_ _2133_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4776_ _2083_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3727_ _1215_ _1221_ _1225_ tree_instances\[16\].u_tree.tree_state\[2\] VGND VGND
+ VPWR VPWR _0017_ sky130_fd_sc_hd__o31a_1
XFILLER_0_99_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6515_ clknet_leaf_2_clk _0298_ net26 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.read_enable
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3658_ _1166_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__clkbuf_1
X_6446_ clknet_leaf_96_clk _0239_ net32 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6377_ clknet_leaf_77_clk _0184_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[1\] sky130_fd_sc_hd__dfrtp_1
X_3589_ _1049_ _1036_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_27_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5328_ _1570_ _2414_ VGND VGND VPWR VPWR _2437_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_179 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5259_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[1\] _1379_ _2399_
+ VGND VGND VPWR VPWR _2401_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_306 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_542 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6766__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkload5_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_66_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_17_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4630_ _1252_ _1989_ _0024_ tree_instances\[19\].u_tree.pipeline_valid\[0\] VGND
+ VGND VPWR VPWR _0192_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_60_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5566__A _2578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6300_ clknet_leaf_14_clk _0109_ net29 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4561_ _1953_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4492_ _1779_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[2\] _1910_
+ _1036_ _1913_ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__a221o_1
X_3512_ tree_instances\[8\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__buf_1
X_6231_ _3113_ VGND VGND VPWR VPWR _3114_ sky130_fd_sc_hd__clkbuf_1
X_3443_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _0973_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6162_ _3070_ VGND VGND VPWR VPWR _3071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3374_ _0911_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
X_5113_ _1451_ _2296_ VGND VGND VPWR VPWR _2303_ sky130_fd_sc_hd__and2_1
X_6093_ _3026_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5044_ _2265_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_88_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6436__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6995_ clknet_leaf_94_clk _0701_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5946_ _2923_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5877_ _2879_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4380__A _1112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4828_ tree_instances\[0\].u_tree.frame_id_in\[0\] VGND VGND VPWR VPWR _2122_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_99_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4759_ tree_instances\[11\].u_tree.frame_id_out\[3\] tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[3\]
+ tree_instances\[11\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2075_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_43_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6429_ clknet_leaf_100_clk _0222_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_491 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4678__A1 _1835_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_14_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_22_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6947__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_72_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3992_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1471_ sky130_fd_sc_hd__inv_2
X_5800_ _2580_ net21 _2583_ VGND VGND VPWR VPWR _2838_ sky130_fd_sc_hd__a21oi_1
X_6780_ clknet_leaf_20_clk _0514_ net25 VGND VGND VPWR VPWR complete_votes\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5731_ tree_instances\[19\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2776_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5662_ complete_votes\[0\] VGND VGND VPWR VPWR _2707_ sky130_fd_sc_hd__inv_2
X_4613_ _1790_ _1937_ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_361 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5593_ _2610_ tree_instances\[13\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2643_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_111_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4544_ tree_instances\[9\].u_tree.tree_state\[1\] tree_instances\[9\].u_tree.tree_state\[2\]
+ _1814_ VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__or3_1
X_4475_ tree_instances\[8\].u_tree.tree_state\[0\] tree_instances\[8\].u_tree.tree_state\[2\]
+ tree_instances\[8\].u_tree.tree_state\[1\] _1897_ VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_40_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6214_ _3103_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6688__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3426_ _0958_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[0\] tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[3\]
+ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__or3_1
X_3357_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _0898_ sky130_fd_sc_hd__buf_1
X_6145_ _3050_ tree_instances\[12\].u_tree.node_data\[12\] _3056_ VGND VGND VPWR VPWR
+ _0643_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6076_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[1\] _1351_ _2989_
+ VGND VGND VPWR VPWR _3017_ sky130_fd_sc_hd__mux2_1
X_5027_ tree_instances\[14\].u_tree.frame_id_out\[1\] tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0735_ VGND VGND VPWR VPWR _2257_ sky130_fd_sc_hd__mux2_1
X_3288_ _0832_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6978_ clknet_leaf_16_clk _0684_ net29 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5929_ tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[3\] _1834_ _0030_ VGND
+ VGND VPWR VPWR _2915_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_106_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_445 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6781__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_537 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4260_ _1728_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
X_3211_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__clkbuf_1
X_4191_ _1662_ VGND VGND VPWR VPWR _1663_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6901_ clknet_leaf_73_clk _0614_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ sky130_fd_sc_hd__dfxtp_1
X_6832_ clknet_leaf_36_clk _0553_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.prediction_out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6959__SET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6763_ clknet_leaf_21_clk _0497_ net24 VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__dfrtp_1
X_3975_ _1436_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__clkbuf_1
X_6694_ clknet_leaf_54_clk _0443_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5714_ _2622_ tree_instances\[18\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2759_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5645_ attack_votes\[0\] VGND VGND VPWR VPWR _2694_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5576_ _2586_ tree_instances\[3\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2626_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4527_ tree_instances\[8\].u_tree.tree_state\[0\] _1034_ tree_instances\[8\].u_tree.tree_state\[1\]
+ VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_111_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4458_ tree_instances\[7\].u_tree.tree_state\[0\] _0969_ VGND VGND VPWR VPWR _1883_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__6451__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3409_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _0944_ sky130_fd_sc_hd__clkbuf_1
X_4389_ _1831_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
X_6128_ _3045_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__clkbuf_1
X_6059_ _2465_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[2\] tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ _2464_ _3001_ VGND VGND VPWR VPWR _3002_ sky130_fd_sc_hd__o221a_1
XFILLER_0_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5781__A2 _2820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_101_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5664__A _2606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3760_ tree_instances\[19\].u_tree.tree_state\[0\] _1251_ _1252_ VGND VGND VPWR VPWR
+ _0065_ sky130_fd_sc_hd__a21o_1
XTAP_TAPCELL_ROW_80_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_27_434 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5430_ _2523_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3691_ _1195_ _0862_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5361_ _2462_ VGND VGND VPWR VPWR _2463_ sky130_fd_sc_hd__clkbuf_1
X_5292_ _2418_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__clkbuf_1
X_4312_ _1778_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4243_ _0845_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4174_ _1645_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_38_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6815_ clknet_leaf_53_clk _0536_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6746_ clknet_leaf_72_clk _0489_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.gen_tree_3.u_tree_rom.node_data\[107\]
+ sky130_fd_sc_hd__dfxtp_1
X_3958_ _1434_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3889_ _1364_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__clkbuf_1
X_6677_ clknet_leaf_63_clk _0427_ net35 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5628_ _2575_ tree_instances\[10\].u_tree.frame_id_out\[0\] _2676_ _2677_ tree_instances\[10\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2678_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_103_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6632__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5559_ _2578_ tree_instances\[20\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2609_
+ sky130_fd_sc_hd__or2b_1
XANTENNA__5279__A1 _2249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_103_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3179__A _0733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_551 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_459 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6373__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6302__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5690__B2 _2659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5690__A1 _2598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4930_ _2111_ VGND VGND VPWR VPWR _2201_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_35_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_164 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_63_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4861_ _2141_ VGND VGND VPWR VPWR _2142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3812_ _1298_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__clkbuf_1
X_6600_ clknet_leaf_60_clk _0364_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4792_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[7\] tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ VGND VGND VPWR VPWR _2095_ sky130_fd_sc_hd__nand2_1
XANTENNA__4953__A0 _1830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6531_ clknet_leaf_31_clk _0038_ net29 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3743_ _0791_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_158 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_554 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6462_ clknet_leaf_100_clk _0250_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.cache_valid
+ sky130_fd_sc_hd__dfxtp_1
X_3674_ _1179_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND
+ VPWR VPWR _1180_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5413_ _2505_ _2506_ _2507_ _2508_ _2509_ VGND VGND VPWR VPWR _2510_ sky130_fd_sc_hd__a221o_1
X_6393_ clknet_leaf_52_clk _0195_ net37 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5344_ state\[1\] VGND VGND VPWR VPWR _2447_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_7_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5275_ tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[1\] _2246_ _0022_ VGND
+ VGND VPWR VPWR _2409_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4226_ _1694_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4157_ _1127_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5681__A1 _2627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4088_ _1562_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__clkbuf_1
Xmax_cap29 net30 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__buf_12
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4383__A _1826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6884__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6813__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6729_ clknet_leaf_67_clk _0477_ net36 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5672__A1 _2714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5672__B2 _2709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_60_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6554__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3390_ _0926_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5060_ _2273_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__clkbuf_1
X_4011_ _1483_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_56 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5962_ tree_instances\[7\].u_tree.pipeline_valid\[0\] tree_instances\[7\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _2931_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4913_ tree_instances\[12\].u_tree.read_enable _2108_ VGND VGND VPWR VPWR _2192_
+ sky130_fd_sc_hd__nand2_4
X_5893_ _2887_ _2889_ _2891_ _2892_ VGND VGND VPWR VPWR _2893_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4844_ _2132_ VGND VGND VPWR VPWR _2133_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_74_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4775_ _1610_ _2030_ VGND VGND VPWR VPWR _2083_ sky130_fd_sc_hd__and2_1
X_3726_ _1224_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6514_ clknet_leaf_99_clk _0297_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.current_node_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6445_ clknet_leaf_23_clk _0238_ net28 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3657_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[5\] _1165_ VGND VGND
+ VPWR VPWR _1166_ sky130_fd_sc_hd__or2_1
X_6376_ clknet_leaf_80_clk _0183_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[0\] sky130_fd_sc_hd__dfrtp_1
X_3588_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1105_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5327_ _2436_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6422__SET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6485__SET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5258_ _2400_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__clkbuf_1
X_5189_ _2362_ VGND VGND VPWR VPWR _2363_ sky130_fd_sc_hd__clkbuf_1
X_4209_ _1648_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND
+ VPWR VPWR _1681_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5709__A2 _2627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_486 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_66_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_109_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_17_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_304 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_69_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6735__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4384__A1 _1827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4560_ _1752_ _1944_ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_404 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_77_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5582__A _2582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4491_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[2\] _1778_ _1774_
+ _1909_ VGND VGND VPWR VPWR _1913_ sky130_fd_sc_hd__a2bb2o_1
X_3511_ _1026_ _1030_ _1033_ tree_instances\[12\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0052_ sky130_fd_sc_hd__a31o_1
X_6230_ _3112_ VGND VGND VPWR VPWR _3113_ sky130_fd_sc_hd__clkbuf_1
X_3442_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _0972_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3373_ _0909_ _0910_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__or2_1
X_6161_ _3069_ VGND VGND VPWR VPWR _3070_ sky130_fd_sc_hd__clkbuf_1
X_5112_ _2302_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5636__A1 _2659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6092_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_data\[107\] tree_instances\[3\].u_tree.u_tree_weight_rom.gen_tree_3.u_tree_rom.node_data\[107\]
+ _3025_ VGND VGND VPWR VPWR _3026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5043_ _1647_ _2222_ VGND VGND VPWR VPWR _2265_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_88_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6994_ clknet_leaf_94_clk _0700_ net27 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6476__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5945_ _1407_ _2553_ VGND VGND VPWR VPWR _2923_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5876_ tree_instances\[1\].u_tree.frame_id_out\[4\] tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[1\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2879_ sky130_fd_sc_hd__mux2_1
XANTENNA__5757__A _2622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6405__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4827_ _2121_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4758_ _2074_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_576 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3709_ tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1209_ sky130_fd_sc_hd__clkbuf_1
X_4689_ _2031_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__clkbuf_1
X_6428_ clknet_leaf_98_clk _0221_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_101_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6359_ clknet_leaf_81_clk _0166_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_42_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_49_Left_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_73_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6987__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_58_Left_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6916__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_11_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3991_ _1469_ _0877_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5730_ _2576_ tree_instances\[19\].u_tree.frame_id_out\[0\] _2772_ _2588_ VGND VGND
+ VPWR VPWR _2775_ sky130_fd_sc_hd__o22a_1
XANTENNA__5577__A _2622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_262 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5661_ _2706_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4612_ _1980_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
X_5592_ current_voting_frame\[4\] tree_instances\[13\].u_tree.frame_id_out\[4\] VGND
+ VGND VPWR VPWR _2642_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4543_ _1000_ _1897_ _1813_ tree_instances\[8\].u_tree.ready_for_next VGND VGND VPWR
+ VPWR _0151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4474_ tree_instances\[8\].u_tree.tree_state\[0\] _0999_ VGND VGND VPWR VPWR _1897_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6213_ tree_instances\[5\].u_tree.frame_id_out\[0\] tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0903_ VGND VGND VPWR VPWR _3103_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3425_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _0958_ sky130_fd_sc_hd__clkbuf_1
X_3356_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _0897_ sky130_fd_sc_hd__clkbuf_1
X_6144_ tree_instances\[12\].u_tree.u_tree_weight_rom.gen_tree_12.u_tree_rom.node_data\[12\]
+ _2112_ _3055_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_data\[12\] VGND
+ VGND VPWR VPWR _3056_ sky130_fd_sc_hd__a22o_1
X_3287_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[5\] tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[4\]
+ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__or2_1
X_6075_ _3016_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__clkbuf_1
X_5026_ _2256_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_92_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_4
X_6977_ clknet_leaf_38_clk _0683_ net29 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5928_ _2914_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5859_ _2869_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_498 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4520__A1 _1835_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6398__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6327__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_83_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_106_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_27_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_55_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_457 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_581 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_387 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_549 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3210_ _0759_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__clkbuf_1
X_4190_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1662_ sky130_fd_sc_hd__inv_2
XANTENNA__6892__SET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6750__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_85_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_74_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_4
X_6900_ clknet_leaf_74_clk _0613_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_106_52 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6831_ clknet_leaf_39_clk _0552_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3974_ _1439_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__clkbuf_1
X_6762_ clknet_leaf_6_clk _0496_ net26 VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_605 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6693_ clknet_leaf_54_clk _0442_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5713_ _2622_ tree_instances\[18\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2758_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_72_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5644_ attack_votes\[0\] attack_votes\[1\] VGND VGND VPWR VPWR _2693_ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_96_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5575_ tree_instances\[3\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2625_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4526_ _1933_ VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4457_ _1882_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3408_ _0936_ _0942_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6838__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4388_ tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[1\] _1830_ _0040_ VGND
+ VGND VPWR VPWR _1831_ sky130_fd_sc_hd__mux2_1
X_6127_ _1344_ _2972_ VGND VGND VPWR VPWR _3045_ sky130_fd_sc_hd__and2_1
X_3339_ _0880_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6255__A1 _1826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6058_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[4\] tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ VGND VGND VPWR VPWR _3001_ sky130_fd_sc_hd__xnor2_1
X_5009_ _2245_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_65_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_24_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_52_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5010__A _1829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_24_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_101_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_51_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3465__A tree_instances\[11\].u_tree.ready_for_next VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4741__A1 _1830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6579__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6508__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_101_Right_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_56_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_4_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_80_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_210 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3690_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5360_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _2462_ sky130_fd_sc_hd__clkbuf_1
X_5291_ tree_instances\[18\].u_tree.frame_id_out\[3\] tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0753_ VGND VGND VPWR VPWR _2418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4311_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1778_ sky130_fd_sc_hd__inv_2
X_4242_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1711_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4173_ _1644_ VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_47_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6814_ clknet_leaf_53_clk _0535_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6745_ clknet_leaf_61_clk _0058_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3957_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_42_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3888_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1371_ sky130_fd_sc_hd__clkbuf_1
X_6676_ clknet_leaf_62_clk _0426_ net35 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5627_ _2582_ tree_instances\[10\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2677_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_257 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5558_ tree_instances\[20\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2608_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_359 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4509_ _1924_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_195 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6672__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire1 clk VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_2
X_5489_ tree_instances\[20\].u_tree.frame_id_out\[4\] tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[20\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2558_ sky130_fd_sc_hd__mux2_1
XANTENNA__6601__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_57_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_1_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_103_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5675__A _2580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_563 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6342__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_69_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_29_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_324 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4860_ _0823_ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_35_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3811_ _1299_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__clkbuf_1
X_6530_ clknet_leaf_30_clk _0037_ net33 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4791_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[7\] tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ VGND VGND VPWR VPWR _2094_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3742_ _1236_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_95 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6461_ clknet_leaf_98_clk _0249_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.pipeline_prediction\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3673_ _1178_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__clkbuf_1
X_5412_ _1481_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[2\] tree_instances\[1\].u_tree.u_tree_weight_rom.cache_valid
+ VGND VGND VPWR VPWR _2509_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6392_ clknet_leaf_96_clk _0194_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.cache_valid
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5343_ _2446_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_99 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5274_ _2408_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__clkbuf_1
X_4225_ _1693_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__clkbuf_1
X_4156_ _1620_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__clkbuf_1
Xmax_cap19 net20 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
X_4087_ _1549_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_108_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4989_ _2233_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__clkbuf_1
X_6728_ clknet_leaf_68_clk _0476_ net36 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_12_Left_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6659_ clknet_leaf_8_clk _0012_ net26 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6853__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5121__A1 _2125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_21_Left_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_60_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_32_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_30_Left_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_12_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6594__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_40_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6523__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4010_ _0867_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5961_ _0755_ _2570_ _1804_ tree_instances\[2\].u_tree.ready_for_next VGND VGND VPWR
+ VPWR _0585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4912_ _2169_ _2191_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_48_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5892_ _1403_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[3\] VGND
+ VGND VPWR VPWR _2892_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4843_ tree_instances\[12\].u_tree.tree_state\[1\] tree_instances\[12\].u_tree.tree_state\[2\]
+ _1810_ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__or3_1
XFILLER_0_28_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4774_ _2082_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3725_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6513_ clknet_leaf_3_clk _0296_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_6444_ clknet_leaf_23_clk _0237_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_9_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3656_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1165_ sky130_fd_sc_hd__buf_1
XFILLER_0_30_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3587_ _1092_ _1097_ _1104_ tree_instances\[9\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0086_ sky130_fd_sc_hd__a31o_1
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6375_ clknet_leaf_19_clk _0182_ net25 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5326_ _1566_ _2414_ VGND VGND VPWR VPWR _2436_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5257_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[0\] _1386_ _2399_
+ VGND VGND VPWR VPWR _2400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4208_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[5\] _1663_ VGND VGND
+ VPWR VPWR _1680_ sky130_fd_sc_hd__nor2_1
X_5188_ _2361_ VGND VGND VPWR VPWR _2362_ sky130_fd_sc_hd__clkbuf_1
X_4139_ _1612_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4394__A _1834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_111_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_load_slew36_A net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_109_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_17_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_316 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_45_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6775__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6704__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3510_ _1031_ _1032_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_77_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4490_ _1774_ _1909_ _1911_ VGND VGND VPWR VPWR _1912_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_25_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3441_ tree_instances\[6\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__clkbuf_1
X_3372_ _0732_ tree_instances\[17\].u_tree.pipeline_valid\[0\] tree_instances\[17\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__o21a_1
X_6160_ tree_instances\[20\].u_tree.read_enable _2894_ VGND VGND VPWR VPWR _3069_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_85_23 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5111_ _1453_ _2296_ VGND VGND VPWR VPWR _2302_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6091_ _2988_ VGND VGND VPWR VPWR _3025_ sky130_fd_sc_hd__clkbuf_1
X_5042_ _2264_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_88_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6993_ clknet_leaf_95_clk _0699_ net32 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5944_ _2922_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5875_ _2878_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_135 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4826_ _1285_ _2070_ VGND VGND VPWR VPWR _2121_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6445__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4757_ tree_instances\[11\].u_tree.frame_id_out\[2\] tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[2\]
+ tree_instances\[11\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3708_ _1007_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__clkbuf_1
X_4688_ tree_instances\[10\].u_tree.frame_id_out\[0\] tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _1136_ VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__mux2_1
X_3639_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1149_ sky130_fd_sc_hd__clkbuf_1
X_6427_ clknet_leaf_96_clk _0220_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6358_ clknet_leaf_80_clk _0165_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[2\]
+ sky130_fd_sc_hd__dfxtp_1
X_5309_ _2426_ VGND VGND VPWR VPWR _2427_ sky130_fd_sc_hd__dlymetal6s2s_1
X_6289_ _3144_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6754__D _0008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_81_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_22_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_72_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3990_ _0868_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6956__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_274 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_466 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5660_ _2705_ _2573_ _2703_ VGND VGND VPWR VPWR _2706_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4611_ _1781_ _1937_ VGND VGND VPWR VPWR _1980_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5593__A _2610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5554__B2 _2603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5591_ _2602_ tree_instances\[13\].u_tree.frame_id_out\[1\] _2639_ _2640_ VGND VGND
+ VPWR VPWR _2641_ sky130_fd_sc_hd__o211a_1
XFILLER_0_111_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4542_ _1943_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5306__A1 _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4473_ tree_instances\[8\].u_tree.tree_state\[1\] tree_instances\[8\].u_tree.current_node_data\[12\]
+ tree_instances\[8\].u_tree.node_data\[12\] _1895_ VGND VGND VPWR VPWR _1896_ sky130_fd_sc_hd__a22o_1
X_6212_ _3004_ _3100_ _3102_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__o21ai_1
X_3424_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3355_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _0896_ sky130_fd_sc_hd__inv_2
X_6143_ _3054_ VGND VGND VPWR VPWR _3055_ sky130_fd_sc_hd__clkbuf_1
X_3286_ _0831_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
X_6074_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[0\] _1325_ _2989_
+ VGND VGND VPWR VPWR _3016_ sky130_fd_sc_hd__mux2_1
X_5025_ tree_instances\[14\].u_tree.frame_id_out\[0\] tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0735_ VGND VGND VPWR VPWR _2256_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5768__A _2610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6697__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6976_ clknet_leaf_81_clk _0682_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cached_data\[107\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6626__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5927_ tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[2\] _2595_ _0030_ VGND
+ VGND VPWR VPWR _2914_ sky130_fd_sc_hd__mux2_1
X_5858_ tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[2\] _2595_ _0026_ VGND
+ VGND VPWR VPWR _2869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5789_ _2821_ _2830_ complete_votes\[3\] net10 VGND VGND VPWR VPWR _2831_ sky130_fd_sc_hd__a2bb2o_1
X_4809_ _2111_ VGND VGND VPWR VPWR _2112_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_17_Right_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_26_Right_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3470__B _0996_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_106_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5678__A _2589_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_27_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6367__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_4_Left_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_116 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_35_Right_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_399 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_44_Right_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6830_ clknet_leaf_40_clk _0551_ net36 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_64 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6761_ clknet_leaf_5_clk _0495_ net26 VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5712_ tree_instances\[18\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2757_ sky130_fd_sc_hd__inv_2
X_3973_ _1452_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_53_Right_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6692_ clknet_leaf_54_clk _0441_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5643_ _2692_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5574_ _2615_ _2618_ _2621_ _2623_ VGND VGND VPWR VPWR _2624_ sky130_fd_sc_hd__and4_1
XTAP_TAPCELL_ROW_96_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_322 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4525_ _1932_ VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__clkbuf_1
X_4456_ _1233_ _1850_ VGND VGND VPWR VPWR _1882_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_62_Right_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3407_ _0941_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__clkbuf_1
X_4387_ _1829_ VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__clkbuf_4
X_3338_ _0878_ _0879_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_293 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6126_ _3044_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6878__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6057_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[7\] _2993_ _2998_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[8\]
+ _2999_ VGND VGND VPWR VPWR _3000_ sky130_fd_sc_hd__o221a_1
X_3269_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__clkbuf_1
X_5008_ tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[0\] _2122_ _0014_ VGND
+ VGND VPWR VPWR _2245_ sky130_fd_sc_hd__mux2_1
XANTENNA__6807__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_77_Left_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_72_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6460__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_71_Right_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5766__B2 _2606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5766__A1 _2619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6959_ clknet_leaf_86_clk _0671_ net30 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_48_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_87_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5945__B _2553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_379 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_631 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_10_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_86_Left_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_80_Right_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_25_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6548__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_4_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_285 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5290_ _2417_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__clkbuf_1
X_4310_ _1041_ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4241_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1710_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_91_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4172_ _1643_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6813_ clknet_leaf_53_clk _0534_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5748__A1 _2576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5748__B2 _2619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3956_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1436_ sky130_fd_sc_hd__clkbuf_1
X_6744_ clknet_leaf_61_clk _0016_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6675_ clknet_leaf_62_clk _0425_ net35 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3887_ _1369_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5626_ tree_instances\[10\].u_tree.frame_id_out\[1\] _2578_ VGND VGND VPWR VPWR _2676_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_5_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5557_ _2598_ tree_instances\[20\].u_tree.frame_id_out\[0\] tree_instances\[20\].u_tree.frame_id_out\[3\]
+ _2606_ VGND VGND VPWR VPWR _2607_ sky130_fd_sc_hd__o22a_1
X_4508_ _1300_ _1840_ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__and2_1
X_5488_ _2557_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4439_ _1868_ _1851_ VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__and2_1
Xwire2 _3007_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
XANTENNA__4397__A tree_instances\[0\].u_tree.frame_id_in\[4\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_111_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6109_ tree_instances\[4\].u_tree.frame_id_out\[0\] tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0849_ VGND VGND VPWR VPWR _3036_ sky130_fd_sc_hd__mux2_1
XANTENNA__6641__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_100 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_103_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_575 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_94_Left_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6729__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6382__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_69_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6311__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3810_ _1293_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4790_ _1711_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[4\] tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ _1691_ _2092_ VGND VGND VPWR VPWR _2093_ sky130_fd_sc_hd__a221o_1
X_3741_ _0792_ _0793_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6460_ clknet_leaf_24_clk _0076_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3672_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1178_ sky130_fd_sc_hd__clkbuf_1
X_5411_ _0878_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[4\] VGND
+ VGND VPWR VPWR _2508_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6391_ clknet_leaf_93_clk _0193_ net25 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_prediction\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5342_ _1018_ _2442_ _2445_ VGND VGND VPWR VPWR _2446_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5273_ tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[0\] _2122_ _0022_ VGND
+ VGND VPWR VPWR _2408_ sky130_fd_sc_hd__mux2_1
X_4224_ _1690_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__clkbuf_1
X_4155_ _1625_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__clkbuf_1
X_4086_ _1560_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5480__B1_N _2553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_108_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4988_ _1679_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[1\] _2231_
+ VGND VGND VPWR VPWR _2233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6727_ clknet_leaf_67_clk _0475_ net36 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3939_ _1408_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6658_ clknet_leaf_1_clk _0011_ net26 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5609_ _2605_ VGND VGND VPWR VPWR _2659_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_103_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6589_ clknet_leaf_83_clk _0042_ net31 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6893__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6822__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_40_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5960_ _2930_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5891_ _1399_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[2\] tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ _1395_ _2890_ VGND VGND VPWR VPWR _2891_ sky130_fd_sc_hd__o221a_1
X_4911_ _2190_ VGND VGND VPWR VPWR _2191_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5596__A _2583_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4842_ tree_instances\[12\].u_tree.tree_state\[0\] _1026_ tree_instances\[12\].u_tree.tree_state\[1\]
+ VGND VGND VPWR VPWR _2131_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_618 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4773_ _1614_ _2030_ VGND VGND VPWR VPWR _2082_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3724_ _0925_ _1222_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__or2_1
X_6512_ clknet_leaf_8_clk _0295_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_6443_ clknet_leaf_23_clk _0236_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3655_ _1163_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3586_ _1100_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__nor2_1
X_6374_ clknet_leaf_15_clk _0181_ net29 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5325_ _2435_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__clkbuf_1
X_5256_ _2362_ VGND VGND VPWR VPWR _2399_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4207_ _1651_ VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5187_ tree_instances\[16\].u_tree.read_enable _2360_ VGND VGND VPWR VPWR _2361_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_97_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4138_ _1611_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__clkbuf_1
X_4069_ _1536_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5953__B _2553_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5878__A0 tree_instances\[1\].u_tree.prediction_out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_111_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6587__SET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_17_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_45_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3440_ tree_instances\[7\].u_tree.tree_state\[0\] _0969_ _0970_ VGND VGND VPWR VPWR
+ _0081_ sky130_fd_sc_hd__a21o_1
XANTENNA__6744__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3371_ tree_instances\[17\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__buf_2
XFILLER_0_0_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5110_ _2301_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__clkbuf_1
X_6090_ _3024_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5041_ _1684_ _2222_ VGND VGND VPWR VPWR _2264_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_51 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6992_ clknet_leaf_96_clk _0698_ net32 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5943_ tree_instances\[2\].u_tree.frame_id_out\[4\] tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[2\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2922_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5874_ tree_instances\[1\].u_tree.frame_id_out\[3\] tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _1227_ VGND VGND VPWR VPWR _2878_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_147 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4825_ _2120_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_478 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_63_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4756_ _2073_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3707_ _1005_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4687_ _2027_ _2028_ _2030_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_43_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3638_ _1143_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_403 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6426_ clknet_leaf_95_clk _0219_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_3_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3569_ _1086_ _1087_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6357_ clknet_leaf_77_clk _0164_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6414__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5308_ tree_instances\[19\].u_tree.tree_state\[1\] tree_instances\[19\].u_tree.tree_state\[2\]
+ _1825_ VGND VGND VPWR VPWR _2426_ sky130_fd_sc_hd__or3_1
X_6288_ _2477_ _3102_ VGND VGND VPWR VPWR _3144_ sky130_fd_sc_hd__and2_1
X_5239_ _2390_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6096__S _0034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_98_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_42_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_504 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_592 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkload3_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_125 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_83_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4610_ _1979_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6996__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6925__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_320 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5590_ current_voting_frame\[0\] tree_instances\[13\].u_tree.frame_id_out\[0\] VGND
+ VGND VPWR VPWR _2640_ sky130_fd_sc_hd__or2b_1
XFILLER_0_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4541_ tree_instances\[8\].u_tree.prediction_out tree_instances\[8\].u_tree.pipeline_prediction\[0\]\[0\]
+ tree_instances\[8\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1943_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4472_ tree_instances\[8\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _1895_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6211_ _3101_ VGND VGND VPWR VPWR _3102_ sky130_fd_sc_hd__clkbuf_2
X_3423_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0956_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5813__S _0004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6142_ _2129_ _2093_ _3051_ _3053_ VGND VGND VPWR VPWR _3054_ sky130_fd_sc_hd__nor4_1
X_3354_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__inv_2
X_6073_ tree_instances\[5\].u_tree.u_tree_weight_rom.gen_tree_5.u_tree_rom.node_data\[107\]
+ _3012_ _3015_ _3013_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__a22o_1
X_3285_ _0829_ _0830_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__or2b_1
X_5024_ _2254_ VGND VGND VPWR VPWR _2255_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6975_ clknet_leaf_83_clk _0681_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[8\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5926_ _2913_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5793__A2 _2820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_242 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5857_ _2868_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5788_ complete_votes\[3\] _2829_ VGND VGND VPWR VPWR _2830_ sky130_fd_sc_hd__xnor2_1
X_4808_ _2110_ VGND VGND VPWR VPWR _2111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4739_ tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[0\] _1827_ _0008_ VGND
+ VGND VPWR VPWR _2064_ sky130_fd_sc_hd__mux2_1
X_6409_ clknet_leaf_10_clk _0211_ net25 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_231 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_128 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_27_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6336__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_105_Left_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_85_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_106_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6760_ clknet_leaf_5_clk _0494_ net26 VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5711_ _2713_ tree_instances\[18\].u_tree.frame_id_out\[1\] tree_instances\[18\].u_tree.frame_id_out\[2\]
+ _2714_ VGND VGND VPWR VPWR _2756_ sky130_fd_sc_hd__a22oi_1
X_3972_ _1446_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__clkbuf_1
X_6691_ clknet_leaf_51_clk _0440_ net35 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5642_ _2597_ attack_votes\[0\] _2691_ VGND VGND VPWR VPWR _2692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_534 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5573_ _2622_ tree_instances\[5\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2623_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_96_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4524_ tree_instances\[8\].u_tree.read_enable VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__inv_2
X_4455_ _1881_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
X_4386_ tree_instances\[0\].u_tree.frame_id_in\[1\] VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__buf_2
X_3406_ _0938_ _0940_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3337_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _0879_ sky130_fd_sc_hd__clkbuf_1
X_6125_ _1347_ _2972_ VGND VGND VPWR VPWR _3044_ sky130_fd_sc_hd__and2_1
XANTENNA__5463__A1 _2122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6056_ _2464_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[5\] tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[0\]
+ _2460_ VGND VGND VPWR VPWR _2999_ sky130_fd_sc_hd__o2bb2a_1
X_3268_ _0811_ _0814_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__nor2_1
X_3199_ _0742_ _0744_ _0750_ _0751_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__o31a_1
X_5007_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_data\[12\] _2191_ _2244_
+ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_348 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6847__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_52_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6958_ clknet_leaf_90_clk _0670_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.prediction_out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5909_ _2163_ _2901_ VGND VGND VPWR VPWR _2905_ sky130_fd_sc_hd__and2_1
X_6889_ clknet_leaf_68_clk _0608_ net36 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.prediction_out
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5518__A2 _1020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6588__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6517__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_297 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4240_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1709_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_91_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5693__A1 _2580_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4171_ _1642_ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__clkbuf_1
X_6812_ clknet_leaf_46_clk _0533_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.cache_valid
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__6940__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3955_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1435_ sky130_fd_sc_hd__clkbuf_1
X_6743_ clknet_leaf_60_clk _0015_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_61 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6674_ clknet_leaf_43_clk _0424_ net35 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3886_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1369_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5625_ _2598_ tree_instances\[10\].u_tree.frame_id_out\[0\] tree_instances\[10\].u_tree.frame_id_out\[1\]
+ _2603_ _2674_ VGND VGND VPWR VPWR _2675_ sky130_fd_sc_hd__a221oi_1
XTAP_TAPCELL_ROW_100_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5556_ _2605_ VGND VGND VPWR VPWR _2606_ sky130_fd_sc_hd__clkbuf_4
X_4507_ _1923_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5487_ tree_instances\[20\].u_tree.frame_id_out\[3\] tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _1197_ VGND VGND VPWR VPWR _2557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4438_ _1867_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__clkbuf_1
X_4369_ _1818_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__inv_2
X_6108_ _3034_ VGND VGND VPWR VPWR _3035_ sky130_fd_sc_hd__dlymetal6s2s_1
X_6039_ _2982_ VGND VGND VPWR VPWR _2983_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_1_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_65_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6681__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_37_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6610__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_144 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_69_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6769__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_178 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6351__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ _1233_ _1234_ _1235_ _0971_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__o31a_1
XFILLER_0_55_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_117 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3671_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1177_ sky130_fd_sc_hd__inv_2
X_5410_ _0877_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[4\] VGND
+ VGND VPWR VPWR _2507_ sky130_fd_sc_hd__or2_1
X_6390_ clknet_leaf_67_clk _0072_ net36 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_93_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5341_ complete_votes\[1\] complete_votes\[3\] _2443_ _2444_ VGND VGND VPWR VPWR
+ _2445_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_71_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5272_ _2407_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5666__A1 _2708_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4223_ _1691_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__clkbuf_1
X_4154_ tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1626_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_86_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4085_ _0743_ VGND VGND VPWR VPWR _1560_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6439__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_62_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5776__B _2820_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_34_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_24_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6726_ clknet_leaf_67_clk _0474_ net36 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4987_ _2232_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3938_ _1417_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__clkbuf_1
X_3869_ _1217_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__inv_2
X_6657_ clknet_leaf_1_clk _0053_ net26 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6588_ clknet_leaf_84_clk _0041_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[8\].u_tree.tree_state\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5608_ _2600_ tree_instances\[8\].u_tree.frame_id_out\[2\] _2656_ _2588_ _2657_ VGND
+ VGND VPWR VPWR _2658_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_39_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5539_ tree_instances\[0\].u_tree.frame_id_in\[0\] tree_instances\[0\].u_tree.frame_id_in\[1\]
+ _2591_ VGND VGND VPWR VPWR _2593_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6862__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_12_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_40_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6532__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5890_ _1396_ _2881_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ _1393_ VGND VGND VPWR VPWR _2890_ sky130_fd_sc_hd__o22a_1
X_4910_ _2189_ VGND VGND VPWR VPWR _2190_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_48_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4841_ _2129_ VGND VGND VPWR VPWR _2130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_31_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4772_ _2081_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__clkbuf_1
X_3723_ _0926_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6511_ clknet_leaf_8_clk _0294_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6442_ clknet_leaf_17_clk _0235_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3654_ _1162_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND
+ VPWR VPWR _1163_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_579 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3585_ _1102_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__clkbuf_1
X_6373_ clknet_leaf_15_clk _0180_ net24 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5324_ _1572_ _2414_ VGND VGND VPWR VPWR _2435_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5255_ _1025_ _2398_ _0044_ tree_instances\[9\].u_tree.pipeline_valid\[0\] VGND VGND
+ VPWR VPWR _0410_ sky130_fd_sc_hd__o2bb2a_1
X_4206_ _1658_ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__clkbuf_1
X_5186_ _2350_ _2352_ _2359_ VGND VGND VPWR VPWR _2360_ sky130_fd_sc_hd__or3b_1
X_4137_ _1602_ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4068_ _1540_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5811__A1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_649 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6709_ clknet_leaf_48_clk _0457_ VGND VGND VPWR VPWR tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[0\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_111_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_111_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_17_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_45_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_77_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_590 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3370_ _0907_ _0729_ _0908_ tree_instances\[4\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0076_ sky130_fd_sc_hd__a31o_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6784__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5040_ _2263_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_88_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6991_ clknet_leaf_82_clk _0697_ net32 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5942_ _2921_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5873_ _2877_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__clkbuf_1
X_4824_ _1286_ _2071_ VGND VGND VPWR VPWR _2120_ sky130_fd_sc_hd__and2_1
XFILLER_0_90_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4755_ tree_instances\[11\].u_tree.frame_id_out\[1\] tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[1\]
+ tree_instances\[11\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2073_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3706_ _1206_ _1100_ _1103_ _1092_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__o31a_1
XFILLER_0_55_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_99_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4686_ _2029_ VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_43_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3637_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__clkbuf_1
X_6425_ clknet_leaf_70_clk _0074_ net36 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3568_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6356_ clknet_leaf_80_clk _0163_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[0\]
+ sky130_fd_sc_hd__dfxtp_1
X_5307_ _2425_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__clkbuf_1
X_3499_ tree_instances\[16\].u_tree.tree_state\[0\] _1022_ _1023_ VGND VGND VPWR VPWR
+ _0059_ sky130_fd_sc_hd__a21o_1
X_6287_ _3143_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__clkbuf_1
X_5238_ _1379_ _2314_ VGND VGND VPWR VPWR _2390_ sky130_fd_sc_hd__and2_1
X_5169_ _2342_ VGND VGND VPWR VPWR _2343_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_95_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_108_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_608 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_129 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_151 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_22_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_18_Left_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_72_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_86_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_71_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_137 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4540_ _1942_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_10_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_4
X_4471_ _1893_ VGND VGND VPWR VPWR _1894_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6965__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_398 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6210_ tree_instances\[5\].u_tree.tree_state\[1\] tree_instances\[5\].u_tree.tree_state\[2\]
+ _1808_ VGND VGND VPWR VPWR _3101_ sky130_fd_sc_hd__or3_1
X_3422_ _0953_ _0954_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__nand2_1
XANTENNA__4514__A1 _1827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6141_ _2099_ _3052_ VGND VGND VPWR VPWR _3053_ sky130_fd_sc_hd__or2b_1
X_3353_ _0887_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__nor2_1
X_6072_ tree_instances\[5\].u_tree.node_data\[107\] tree_instances\[5\].u_tree.u_tree_weight_rom.cached_data\[107\]
+ _3014_ VGND VGND VPWR VPWR _3015_ sky130_fd_sc_hd__mux2_1
X_3284_ _0731_ tree_instances\[12\].u_tree.pipeline_valid\[0\] tree_instances\[12\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5023_ tree_instances\[14\].u_tree.tree_state\[1\] tree_instances\[14\].u_tree.tree_state\[2\]
+ _1817_ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_77_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6974_ clknet_leaf_94_clk _0680_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_5925_ tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[1\] _1829_ _0030_ VGND
+ VGND VPWR VPWR _2913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5856_ tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[1\] _1829_ _0026_ VGND
+ VGND VPWR VPWR _2868_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4807_ _2109_ VGND VGND VPWR VPWR _2110_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_3_Right_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5787_ _2823_ _2444_ VGND VGND VPWR VPWR _2829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4738_ _2063_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4669_ _2019_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_346 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6408_ clknet_leaf_91_clk _0210_ net25 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6635__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6339_ clknet_leaf_90_clk _0147_ net31 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_68_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_94_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_55_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_301 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3495__A _1020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_313 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6376__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6305__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_19 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6739__SET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_59_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_85_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3971_ _1448_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5710_ _2748_ _2754_ _2652_ _2679_ VGND VGND VPWR VPWR _2755_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6690_ clknet_leaf_51_clk _0439_ net35 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5641_ _1018_ _2690_ VGND VGND VPWR VPWR _2691_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_546 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5572_ current_voting_frame\[0\] VGND VGND VPWR VPWR _2622_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_96_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4523_ _1931_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
X_4454_ _1880_ _1850_ VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__and2_1
X_4385_ _1828_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
X_3405_ _0939_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__clkbuf_1
X_3336_ _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__clkbuf_1
X_6124_ _3043_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__clkbuf_1
X_6055_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[8\] VGND VGND VPWR
+ VPWR _2998_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5006_ _2241_ tree_instances\[13\].u_tree.u_tree_weight_rom.gen_tree_13.u_tree_rom.node_data\[12\]
+ _2243_ VGND VGND VPWR VPWR _2244_ sky130_fd_sc_hd__and3_1
X_3267_ _0813_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__clkbuf_1
X_3198_ tree_instances\[18\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6957_ clknet_leaf_87_clk _0669_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_52_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6888_ clknet_leaf_89_clk _0607_ net30 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5908_ _2904_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__clkbuf_1
X_5839_ _2859_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6887__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6816__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_4_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_80_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_80_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6557__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4170_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1642_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_91_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6811_ clknet_leaf_35_clk _0532_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_prediction\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3954_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1434_ sky130_fd_sc_hd__clkbuf_1
X_6742_ clknet_leaf_60_clk _0057_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
X_3885_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1368_ sky130_fd_sc_hd__inv_2
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6673_ clknet_leaf_62_clk _0423_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6980__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5624_ _2610_ tree_instances\[10\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2674_
+ sky130_fd_sc_hd__xor2_1
XTAP_TAPCELL_ROW_100_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5555_ current_voting_frame\[3\] VGND VGND VPWR VPWR _2605_ sky130_fd_sc_hd__inv_2
X_4506_ _1305_ _1840_ VGND VGND VPWR VPWR _1923_ sky130_fd_sc_hd__and2_1
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5486_ _2556_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__clkbuf_1
X_4437_ _1866_ VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__clkbuf_1
X_4368_ _1112_ tree_instances\[0\].u_tree.pipeline_valid\[0\] tree_instances\[0\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__or3b_2
X_6107_ tree_instances\[4\].u_tree.tree_state\[1\] tree_instances\[4\].u_tree.tree_state\[2\]
+ _1807_ VGND VGND VPWR VPWR _3034_ sky130_fd_sc_hd__or3_1
XANTENNA__3695__A1 _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3319_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _0862_ sky130_fd_sc_hd__buf_1
X_4299_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[0\] tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[2\]
+ VGND VGND VPWR VPWR _1766_ sky130_fd_sc_hd__nand2b_1
X_6038_ _2968_ _2947_ VGND VGND VPWR VPWR _2982_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_1_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_224 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_340 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_9_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_69_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6738__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3670_ _1175_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__buf_1
XANTENNA__6391__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6320__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5340_ complete_votes\[0\] complete_votes\[2\] VGND VGND VPWR VPWR _2444_ sky130_fd_sc_hd__nand2_1
X_5271_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[7\] _1376_ _2399_
+ VGND VGND VPWR VPWR _2407_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4222_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1691_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4153_ _1125_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__clkbuf_1
X_4084_ _1558_ VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_62_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4986_ _1666_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[0\] _2231_
+ VGND VGND VPWR VPWR _2232_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_34_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6479__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6725_ clknet_leaf_35_clk _0473_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3937_ _1392_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6408__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6656_ clknet_leaf_19_clk _0410_ net24 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3868_ _1343_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_46_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3799_ tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_430 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6587_ clknet_leaf_84_clk _0083_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[8\].u_tree.tree_state\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_33_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5607_ _2578_ tree_instances\[8\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2657_
+ sky130_fd_sc_hd__xor2_1
X_5538_ _1827_ _2591_ _1830_ VGND VGND VPWR VPWR _2592_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_181 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5469_ tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[3\] _2249_ _0028_ VGND
+ VGND VPWR VPWR _2546_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_6_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6831__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_75_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4856__A0 tree_instances\[12\].u_tree.prediction_out VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XANTENNA__6919__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_48_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4840_ tree_instances\[12\].u_tree.read_enable VGND VGND VPWR VPWR _2129_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6572__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_31_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5584__A1 _2627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6501__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4771_ _1608_ _2030_ VGND VGND VPWR VPWR _2081_ sky130_fd_sc_hd__and2_1
X_6510_ clknet_leaf_8_clk _0293_ net27 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3722_ _1218_ _1220_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6441_ clknet_leaf_23_clk _0234_ net24 VGND VGND VPWR VPWR tree_instances\[11\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3653_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1162_ sky130_fd_sc_hd__clkbuf_1
X_6372_ clknet_leaf_15_clk _0179_ net29 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5323_ _2434_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__clkbuf_1
X_3584_ _1101_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5254_ tree_instances\[9\].u_tree.pipeline_valid\[0\] tree_instances\[9\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _2398_ sky130_fd_sc_hd__nand2_1
X_5185_ tree_instances\[16\].u_tree.u_tree_weight_rom.cache_valid _2356_ _2358_ VGND
+ VGND VPWR VPWR _2359_ sky130_fd_sc_hd__and3_1
X_4205_ _1655_ VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__clkbuf_1
X_4136_ _1600_ VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__clkbuf_1
X_4067_ _1541_ VGND VGND VPWR VPWR _1543_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire20 _2661_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_522 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4969_ tree_instances\[13\].u_tree.frame_id_out\[0\] tree_instances\[13\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _1114_ VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__mux2_1
X_6708_ clknet_leaf_74_clk _0456_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.u_tree_weight_rom.cache_valid
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_46_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6639_ clknet_leaf_41_clk _0398_ net36 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_111_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_110_Right_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_17_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_70_clk_A clknet_3_5__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_45_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_85_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_107_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_23_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6753__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6990_ clknet_leaf_96_clk _0696_ net32 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_38_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5941_ tree_instances\[2\].u_tree.frame_id_out\[3\] tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0755_ VGND VGND VPWR VPWR _2921_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_606 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5872_ tree_instances\[1\].u_tree.frame_id_out\[2\] tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _1227_ VGND VGND VPWR VPWR _2877_ sky130_fd_sc_hd__mux2_1
X_4823_ _2119_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5557__B2 _2606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5557__A1 _2598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4754_ _2072_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3705_ _1093_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND
+ VPWR VPWR _1206_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_99_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4685_ tree_instances\[10\].u_tree.tree_state\[1\] tree_instances\[10\].u_tree.tree_state\[2\]
+ _1819_ VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__or3_1
X_3636_ _1144_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__or2_1
X_6424_ clknet_leaf_71_clk _0032_ net38 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3567_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1086_ sky130_fd_sc_hd__clkbuf_1
X_6355_ clknet_leaf_30_clk _0162_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5306_ tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[4\] _2251_ _0024_ VGND
+ VGND VPWR VPWR _2425_ sky130_fd_sc_hd__mux2_1
X_6286_ _2490_ _3102_ VGND VGND VPWR VPWR _3143_ sky130_fd_sc_hd__and2_1
X_5237_ _2389_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__clkbuf_1
X_3498_ tree_instances\[16\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__buf_2
X_5168_ _2341_ VGND VGND VPWR VPWR _2342_ sky130_fd_sc_hd__clkbuf_1
X_5099_ _2295_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5798__A _2713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4119_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1594_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6423__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_42_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3468__D tree_instances\[16\].u_tree.ready_for_next VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_42_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_22_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5720__B2 _2709_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_load_slew34_A net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_83_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_149 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4470_ _1892_ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5711__A1 _2713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5711__B2 _2714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3421_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[5\] tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[6\]
+ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3352_ _0889_ _0892_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__nand2_1
X_6140_ tree_instances\[12\].u_tree.u_tree_weight_rom.cache_valid _2100_ _2101_ _2102_
+ VGND VGND VPWR VPWR _3052_ sky130_fd_sc_hd__and4_1
XFILLER_0_0_433 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6071_ tree_instances\[5\].u_tree.read_enable VGND VGND VPWR VPWR _3014_ sky130_fd_sc_hd__clkbuf_1
X_3283_ tree_instances\[12\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__buf_2
X_5022_ _2253_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_73 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6973_ clknet_leaf_94_clk _0679_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_5924_ _2912_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5855_ _2867_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4806_ tree_instances\[12\].u_tree.read_enable _2108_ VGND VGND VPWR VPWR _2109_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5786_ _2828_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4737_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_data\[12\] tree_instances\[10\].u_tree.u_tree_weight_rom.gen_tree_10.u_tree_rom.node_data\[12\]
+ _2054_ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4668_ _1636_ _2012_ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__and2_1
XANTENNA__6384__SET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3619_ _1128_ _1132_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6407_ clknet_leaf_91_clk _0209_ net25 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4599_ tree_instances\[8\].u_tree.current_node_data\[12\] tree_instances\[8\].u_tree.node_data\[12\]
+ _1034_ VGND VGND VPWR VPWR _1974_ sky130_fd_sc_hd__mux2_1
X_6338_ clknet_leaf_90_clk _0146_ net31 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6269_ _3134_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6675__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6604__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5769__A1 _2575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5769__B2 _2600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6345__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_13_Right_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4680__A1 _1837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_34 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_85_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3970_ _1447_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_586 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5640_ _2614_ _2636_ net11 VGND VGND VPWR VPWR _2690_ sky130_fd_sc_hd__or3b_1
XFILLER_0_53_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_22_Right_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_75 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5571_ _2619_ tree_instances\[5\].u_tree.frame_id_out\[2\] _2620_ VGND VGND VPWR
+ VPWR _2621_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_96_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4522_ tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[4\] _1837_ _0042_ VGND
+ VGND VPWR VPWR _1931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4453_ _1879_ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6457__SET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3404_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0939_ sky130_fd_sc_hd__buf_1
XFILLER_0_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4384_ tree_instances\[7\].u_tree.pipeline_frame_id\[0\]\[0\] _1827_ _0040_ VGND
+ VGND VPWR VPWR _1828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3335_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _0877_ sky130_fd_sc_hd__buf_1
X_6123_ _1350_ _2972_ VGND VGND VPWR VPWR _3043_ sky130_fd_sc_hd__and2_1
XPHY_EDGE_ROW_0_Left_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6054_ _1247_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[6\] tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[8\]
+ _2472_ VGND VGND VPWR VPWR _2997_ sky130_fd_sc_hd__o22a_1
XPHY_EDGE_ROW_31_Right_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3266_ _0812_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_37_Left_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_72 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5005_ _2242_ VGND VGND VPWR VPWR _2243_ sky130_fd_sc_hd__clkbuf_1
X_3197_ _0749_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6956_ clknet_leaf_87_clk _0668_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[5\].u_tree.frame_id_out\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_52_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5907_ _2161_ _2901_ VGND VGND VPWR VPWR _2904_ sky130_fd_sc_hd__and2_1
X_6887_ clknet_leaf_13_clk _0606_ net30 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5838_ _1527_ _2427_ VGND VGND VPWR VPWR _2859_ sky130_fd_sc_hd__and2_1
XFILLER_0_91_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_40_Right_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_46_Left_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5769_ _2575_ tree_instances\[7\].u_tree.frame_id_out\[0\] tree_instances\[7\].u_tree.frame_id_out\[2\]
+ _2600_ _2813_ VGND VGND VPWR VPWR _2814_ sky130_fd_sc_hd__o221a_1
XANTENNA__5923__A1 _1826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_385 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_16_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_17_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6856__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_EDGE_ROW_55_Left_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5035__B _2222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6100__A1 _1834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6792__D _0004_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_4_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_64_Left_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_394 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_54_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_483 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6597__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_73_Left_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6526__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_82_Left_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6810_ clknet_leaf_79_clk _0531_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
X_6741_ clknet_leaf_35_clk _0488_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3953_ _1419_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__clkbuf_1
X_3884_ _1216_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__buf_1
X_6672_ clknet_leaf_62_clk _0422_ net35 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5623_ _2585_ tree_instances\[10\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2673_
+ sky130_fd_sc_hd__xnor2_1
XTAP_TAPCELL_ROW_100_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_14_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5554_ _2600_ tree_instances\[20\].u_tree.frame_id_out\[2\] tree_instances\[20\].u_tree.frame_id_out\[1\]
+ _2603_ VGND VGND VPWR VPWR _2604_ sky130_fd_sc_hd__o2bb2a_1
X_4505_ _1922_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5485_ tree_instances\[20\].u_tree.frame_id_out\[2\] tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _1197_ VGND VGND VPWR VPWR _2556_ sky130_fd_sc_hd__mux2_1
X_4436_ _1865_ VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_41 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4367_ _1817_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3318_ _0857_ _0860_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__nor2_1
X_6106_ _3033_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__clkbuf_1
X_4298_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1765_ sky130_fd_sc_hd__clkbuf_1
X_6037_ _2873_ tree_instances\[1\].u_tree.node_data\[12\] tree_instances\[1\].u_tree.u_tree_weight_rom.cached_data\[12\]
+ _2981_ _2532_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__a221o_1
X_3249_ _0789_ _0797_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_37_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6939_ clknet_leaf_26_clk _0651_ net24 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_353 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6690__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_69_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6778__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6707__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_93_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5270_ _2406_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4221_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1690_ sky130_fd_sc_hd__clkbuf_1
X_4152_ _1131_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_30 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4083_ _0746_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_90_Left_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4985_ _2189_ VGND VGND VPWR VPWR _2231_ sky130_fd_sc_hd__clkbuf_2
XTAP_TAPCELL_ROW_34_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6724_ clknet_leaf_35_clk _0472_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3936_ _1397_ _1409_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6655_ clknet_leaf_37_clk _0060_ net30 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3867_ _1330_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6586_ clknet_leaf_65_clk _0093_ net36 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6448__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_152 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3798_ _1287_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
X_5606_ tree_instances\[8\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2656_ sky130_fd_sc_hd__inv_2
X_5537_ _1827_ _2591_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__xor2_1
XFILLER_0_14_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5468_ _2545_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4419_ _1852_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5399_ tree_instances\[20\].u_tree.tree_state\[1\] tree_instances\[20\].u_tree.current_node_data\[12\]
+ tree_instances\[20\].u_tree.node_data\[12\] _2497_ VGND VGND VPWR VPWR _2498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6800__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_239 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_75_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5281__A1 _2251_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4770_ _2080_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_31_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3721_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[3\] _1219_ VGND VGND
+ VPWR VPWR _1220_ sky130_fd_sc_hd__nor2_1
XFILLER_0_99_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3652_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__clkbuf_1
X_6440_ clknet_leaf_93_clk _0233_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.current_node_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3583_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[5\] tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[4\]
+ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__or2_1
X_6371_ clknet_leaf_15_clk _0178_ net29 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_11_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5322_ _1571_ _2414_ VGND VGND VPWR VPWR _2434_ sky130_fd_sc_hd__and2_1
XFILLER_0_51_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5253_ _0909_ _2397_ _2365_ tree_instances\[17\].u_tree.ready_for_next VGND VGND
+ VPWR VPWR _0409_ sky130_fd_sc_hd__a22o_1
X_5184_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[6\] _2347_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ _1368_ _2357_ VGND VGND VPWR VPWR _2358_ sky130_fd_sc_hd__o221a_1
X_4204_ _1675_ VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4135_ _1601_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__clkbuf_1
X_4066_ _1538_ VGND VGND VPWR VPWR _1542_ sky130_fd_sc_hd__clkbuf_1
Xwire10 _2728_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_78_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6629__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4968_ _2219_ _2220_ _2222_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__o21ai_1
X_3919_ _1398_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__inv_2
X_4899_ _0963_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[4\] VGND
+ VGND VPWR VPWR _2179_ sky130_fd_sc_hd__nor2_1
X_6707_ clknet_leaf_69_clk _0455_ net38 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_prediction\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_3_2__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6638_ clknet_leaf_64_clk _0397_ net35 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6569_ clknet_leaf_61_clk _0338_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4838__A1 _1837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5043__B _2222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_69_Right_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_77_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_78_Right_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4829__A1 _2122_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_10 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5940_ _2920_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_87_Right_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_618 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6793__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5871_ _2876_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6722__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4822_ _1281_ _2071_ VGND VGND VPWR VPWR _2119_ sky130_fd_sc_hd__and2_1
X_4753_ tree_instances\[11\].u_tree.frame_id_out\[0\] tree_instances\[11\].u_tree.pipeline_frame_id\[0\]\[0\]
+ tree_instances\[11\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3704_ _1200_ _1147_ _1204_ _1205_ _1140_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__o41a_1
XANTENNA__6004__S _0032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_99_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6423_ clknet_leaf_71_clk _0031_ net38 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4684_ tree_instances\[10\].u_tree.tree_state\[0\] _1172_ tree_instances\[10\].u_tree.tree_state\[1\]
+ VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__o21ba_1
X_3635_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1145_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_96_Right_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3566_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6354_ clknet_leaf_100_clk _0161_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.gen_tree_12.u_tree_rom.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_24_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3497_ _0732_ tree_instances\[16\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _1022_ sky130_fd_sc_hd__or2_1
X_5305_ _2424_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6285_ _3142_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__clkbuf_1
X_5236_ _1386_ _2314_ VGND VGND VPWR VPWR _2389_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5493__B2 tree_instances\[20\].u_tree.ready_for_next VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
X_5167_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _2341_ sky130_fd_sc_hd__clkbuf_1
X_5098_ tree_instances\[16\].u_tree.u_tree_weight_rom.cache_valid tree_instances\[16\].u_tree.read_enable
+ VGND VGND VPWR VPWR _2295_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4118_ _1592_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__clkbuf_1
X_4049_ _1520_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_42_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6463__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_267 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_100_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_72_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_83_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3420_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _0953_ sky130_fd_sc_hd__inv_2
X_3351_ _0890_ _0891_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6070_ _3005_ VGND VGND VPWR VPWR _3013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3282_ _0802_ _0809_ _0828_ tree_instances\[2\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0072_ sky130_fd_sc_hd__a31o_1
X_5021_ tree_instances\[13\].u_tree.current_node_data\[12\] tree_instances\[13\].u_tree.node_data\[12\]
+ _0968_ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6972_ clknet_leaf_95_clk _0678_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_45_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5923_ tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[0\] _1826_ _0030_ VGND
+ VGND VPWR VPWR _2912_ sky130_fd_sc_hd__mux2_1
X_5854_ tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[0\] _1826_ _0026_ VGND
+ VGND VPWR VPWR _2867_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_48_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4805_ _2093_ _2099_ _2103_ _2107_ VGND VGND VPWR VPWR _2108_ sky130_fd_sc_hd__or4bb_2
X_5785_ _2827_ _2826_ _2825_ VGND VGND VPWR VPWR _2828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4736_ _2062_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__clkbuf_1
X_4667_ _2018_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3618_ _1129_ _1131_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__nor2_1
X_6406_ clknet_leaf_93_clk _0208_ net26 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.read_enable
+ sky130_fd_sc_hd__dfrtp_1
X_4598_ _1973_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
X_6337_ clknet_leaf_90_clk _0145_ net31 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3549_ _1068_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6268_ tree_instances\[6\].u_tree.frame_id_out\[0\] tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0932_ VGND VGND VPWR VPWR _3134_ sky130_fd_sc_hd__mux2_1
X_5219_ _2380_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__clkbuf_1
X_6199_ tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[0\] _1826_ _0036_ VGND
+ VGND VPWR VPWR _3095_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_84_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5218__A1 _2125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6644__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_55_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_99_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_520 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_37_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_85_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6385__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkload1_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_106_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6314__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4968__B1 _2222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5570_ _2585_ tree_instances\[5\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2620_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_25_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4521_ _1930_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_96_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4452_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1879_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3403_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4383_ _1826_ VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3334_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _0876_ sky130_fd_sc_hd__clkbuf_1
X_6122_ _3042_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__clkbuf_1
X_6053_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND VGND VPWR
+ VPWR _2996_ sky130_fd_sc_hd__inv_2
X_3265_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _0812_ sky130_fd_sc_hd__clkbuf_1
X_5004_ _2188_ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__clkbuf_1
X_3196_ _0748_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4959__A0 _1837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6955_ clknet_leaf_87_clk _0667_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[5\].u_tree.frame_id_out\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_52_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5906_ _2903_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5620__B2 _2582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6886_ clknet_leaf_89_clk _0605_ net29 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_EDGE_ROW_101_Left_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5837_ _2530_ _2531_ tree_instances\[1\].u_tree.u_tree_weight_rom.cache_valid VGND
+ VGND VPWR VPWR _0533_ sky130_fd_sc_hd__a21o_1
XFILLER_0_91_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5768_ _2610_ tree_instances\[7\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2813_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_397 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4719_ _2049_ VGND VGND VPWR VPWR _2053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5699_ _2659_ tree_instances\[17\].u_tree.frame_id_out\[3\] _2742_ _2743_ tree_instances\[17\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2744_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_32_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_110_Left_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6825__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_646 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_4_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_105_Right_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5611__A1 _2631_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_133 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_80_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6102__S _0034_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_91_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6566__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6740_ clknet_leaf_68_clk _0099_ net36 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_362 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3952_ _1415_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3883_ _1365_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__clkbuf_1
X_6671_ clknet_leaf_62_clk _0421_ net37 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5622_ tree_instances\[8\].u_tree.prediction_out _2654_ net20 _2671_ tree_instances\[12\].u_tree.prediction_out
+ VGND VGND VPWR VPWR _2672_ sky130_fd_sc_hd__a32o_1
XTAP_TAPCELL_ROW_100_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5553_ _2602_ VGND VGND VPWR VPWR _2603_ sky130_fd_sc_hd__clkbuf_4
X_4504_ _1309_ _1840_ VGND VGND VPWR VPWR _1922_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6012__S _0032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5484_ _2555_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__clkbuf_1
X_4435_ _0973_ VGND VGND VPWR VPWR _1865_ sky130_fd_sc_hd__clkbuf_1
X_4366_ _1112_ tree_instances\[14\].u_tree.pipeline_valid\[0\] tree_instances\[14\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__or3b_2
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3317_ _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__clkbuf_1
X_6105_ tree_instances\[3\].u_tree.current_node_data\[107\] tree_instances\[3\].u_tree.node_data\[107\]
+ _3032_ VGND VGND VPWR VPWR _3033_ sky130_fd_sc_hd__mux2_1
XANTENNA__6094__A1 _1826_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4297_ _1763_ VGND VGND VPWR VPWR _1764_ sky130_fd_sc_hd__clkbuf_1
X_6036_ _2980_ VGND VGND VPWR VPWR _2981_ sky130_fd_sc_hd__clkbuf_1
X_3248_ _0791_ _0796_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__nand2_1
XFILLER_0_96_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3179_ _0733_ tree_instances\[14\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _0734_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_1_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6938_ clknet_leaf_26_clk _0650_ net24 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6869_ clknet_leaf_73_clk _0588_ VGND VGND VPWR VPWR tree_instances\[3\].u_tree.u_tree_weight_rom.cache_valid
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_183 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_9_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_4_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_421 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_307 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_373 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4220_ _1689_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_4151_ _1622_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4082_ _1556_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_102_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4984_ _1822_ _1114_ _2230_ tree_instances\[13\].u_tree.pipeline_valid\[0\] VGND
+ VGND VPWR VPWR _0306_ sky130_fd_sc_hd__o2bb2a_1
XTAP_TAPCELL_ROW_34_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6723_ clknet_leaf_34_clk _0471_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_62_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3935_ _1414_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6654_ clknet_leaf_37_clk _0018_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3866_ _1338_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__clkbuf_1
X_5605_ _2575_ tree_instances\[8\].u_tree.frame_id_out\[0\] tree_instances\[8\].u_tree.frame_id_out\[3\]
+ _2605_ VGND VGND VPWR VPWR _2655_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6585_ clknet_leaf_61_clk _0354_ net38 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3797_ tree_instances\[8\].u_tree.prediction_valid _1000_ VGND VGND VPWR VPWR _1287_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5536_ state\[1\] _2441_ VGND VGND VPWR VPWR _2591_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_60 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5467_ tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[2\] _2125_ _0028_ VGND
+ VGND VPWR VPWR _2545_ sky130_fd_sc_hd__mux2_1
X_4418_ _1849_ _1851_ VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__and2_1
XANTENNA__6488__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6417__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_6_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5398_ _0756_ VGND VGND VPWR VPWR _2497_ sky130_fd_sc_hd__clkbuf_1
X_4349_ _1808_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__inv_2
X_6019_ _2971_ VGND VGND VPWR VPWR _2972_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_424 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6840__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_102_172 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_251 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5520__A _2578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_284 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3720_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1219_ sky130_fd_sc_hd__buf_1
XFILLER_0_83_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_40_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_28_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3651_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[3\] _1159_ VGND VGND
+ VPWR VPWR _1160_ sky130_fd_sc_hd__or2_1
X_3582_ _1098_ _1099_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_11_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6370_ clknet_leaf_84_clk _0177_ net39 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.current_node_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_5321_ _2433_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6581__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_109 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5252_ _0910_ VGND VGND VPWR VPWR _2397_ sky130_fd_sc_hd__inv_2
XANTENNA__6510__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5183_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[4\] tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ VGND VGND VPWR VPWR _2357_ sky130_fd_sc_hd__xnor2_1
X_4203_ _1674_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4134_ _1587_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4745__S _0008_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4065_ _1533_ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__clkbuf_1
Xwire11 net12 VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_1
Xwire22 net23 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_78_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_19_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_93_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4967_ _2221_ VGND VGND VPWR VPWR _2222_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_46_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_31_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_4
X_3918_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1398_ sky130_fd_sc_hd__clkbuf_1
X_6706_ clknet_leaf_91_clk _0454_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_4898_ _1640_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[5\] VGND
+ VGND VPWR VPWR _2178_ sky130_fd_sc_hd__and2_1
X_6637_ clknet_leaf_64_clk _0396_ net35 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3849_ _1333_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_437 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6669__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_357 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6568_ clknet_leaf_67_clk _0337_ net36 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5519_ current_voting_frame\[1\] VGND VGND VPWR VPWR _2578_ sky130_fd_sc_hd__clkbuf_4
X_6499_ clknet_leaf_100_clk _0282_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.cached_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_14_295 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_98_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_276 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_22_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_77_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6339__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_89_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_88_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_88_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5870_ tree_instances\[1\].u_tree.frame_id_out\[1\] tree_instances\[1\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _1227_ VGND VGND VPWR VPWR _2876_ sky130_fd_sc_hd__mux2_1
X_4821_ _2118_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_16_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6203__A1 _2595_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4752_ _2070_ VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__dlymetal6s2s_1
Xclkbuf_leaf_13_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_42 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_237 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3703_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[1\] tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[2\]
+ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4683_ _2026_ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_99_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3634_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1144_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6762__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6422_ clknet_leaf_71_clk _0073_ net38 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_50_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3565_ _1082_ _1083_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6353_ clknet_leaf_70_clk _0160_ net38 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5304_ tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[3\] _2249_ _0024_ VGND
+ VGND VPWR VPWR _2424_ sky130_fd_sc_hd__mux2_1
X_3496_ _1021_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__buf_2
X_6284_ _2468_ _3102_ VGND VGND VPWR VPWR _3142_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_110_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5235_ _2388_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_287 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5166_ _2339_ VGND VGND VPWR VPWR _2340_ sky130_fd_sc_hd__clkbuf_1
X_5097_ _2294_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4117_ _1577_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__clkbuf_1
X_4048_ _1524_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5999_ _2895_ VGND VGND VPWR VPWR _2959_ sky130_fd_sc_hd__buf_1
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_22_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_22_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_83_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4747__A1 _1837_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_508 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3350_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0891_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5020_ _2252_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3281_ _0820_ _0827_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_2_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6971_ clknet_leaf_96_clk _0677_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ sky130_fd_sc_hd__dfxtp_1
X_5922_ _2911_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5853_ _2866_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_513 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6943__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5784_ _2826_ _0000_ VGND VGND VPWR VPWR _2827_ sky130_fd_sc_hd__nor2_1
X_4804_ tree_instances\[12\].u_tree.u_tree_weight_rom.cache_valid _2104_ _2105_ _2106_
+ VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_557 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4735_ _1604_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[7\] _2009_
+ VGND VGND VPWR VPWR _2062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4666_ _1623_ _2012_ VGND VGND VPWR VPWR _2018_ sky130_fd_sc_hd__and2_1
X_3617_ _1130_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__clkbuf_1
X_4597_ tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[4\] _1837_ _0044_ VGND
+ VGND VPWR VPWR _1973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6405_ clknet_leaf_91_clk _0207_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3548_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6336_ clknet_leaf_79_clk _0144_ net39 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.read_enable
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3479_ tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1006_ sky130_fd_sc_hd__clkbuf_1
X_6267_ _3133_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__clkbuf_1
X_6198_ _3094_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__clkbuf_1
X_5218_ tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[2\] _2125_ _0020_ VGND
+ VGND VPWR VPWR _2380_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5149_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _2323_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6684__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_35_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_85_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_600 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_260 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4520_ tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[3\] _1835_ _0042_ VGND
+ VGND VPWR VPWR _1930_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_96_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4451_ _1878_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3402_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _0937_ sky130_fd_sc_hd__buf_1
XFILLER_0_40_157 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4382_ tree_instances\[0\].u_tree.frame_id_in\[0\] VGND VGND VPWR VPWR _1826_ sky130_fd_sc_hd__clkbuf_4
X_6121_ _1351_ _2972_ VGND VGND VPWR VPWR _3042_ sky130_fd_sc_hd__and2_1
X_3333_ _0874_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6052_ _2450_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[1\] tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[2\]
+ _2465_ _2994_ VGND VGND VPWR VPWR _2995_ sky130_fd_sc_hd__a221oi_1
XPHY_EDGE_ROW_7_Right_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3264_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__clkbuf_1
X_5003_ _2240_ VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__clkbuf_1
X_3195_ _0745_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6954_ clknet_leaf_88_clk _0666_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[5\].u_tree.frame_id_out\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_105_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_24_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5905_ _2149_ _2901_ VGND VGND VPWR VPWR _2903_ sky130_fd_sc_hd__and2_1
X_6885_ clknet_leaf_12_clk _0604_ net29 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_52_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5836_ _2858_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5767_ _2709_ tree_instances\[7\].u_tree.frame_id_out\[3\] _2811_ VGND VGND VPWR
+ VPWR _2812_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5698_ _2588_ tree_instances\[17\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2743_
+ sky130_fd_sc_hd__xnor2_1
X_4718_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_data\[12\] _2048_ _2052_
+ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a21o_1
XFILLER_0_102_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4649_ _1165_ _1999_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ _1595_ _2006_ VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_81 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6319_ clknet_leaf_14_clk _0105_ net29 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5613__A _2610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_4_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_80_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4838__S _0010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_91_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3951_ _0767_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3882_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_374 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_73_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6670_ clknet_leaf_63_clk _0420_ net35 VGND VGND VPWR VPWR tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5621_ _2664_ _2667_ _2670_ VGND VGND VPWR VPWR _2671_ sky130_fd_sc_hd__and3_1
XTAP_TAPCELL_ROW_100_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5552_ current_voting_frame\[1\] VGND VGND VPWR VPWR _2602_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4503_ _1921_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_83_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5483_ tree_instances\[20\].u_tree.frame_id_out\[1\] tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _1197_ VGND VGND VPWR VPWR _2555_ sky130_fd_sc_hd__mux2_1
X_4434_ _1864_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4365_ _1816_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3316_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[0\] _0858_ VGND VGND
+ VPWR VPWR _0859_ sky130_fd_sc_hd__or2_1
X_6104_ _2932_ VGND VGND VPWR VPWR _3032_ sky130_fd_sc_hd__clkbuf_1
X_6035_ _2979_ VGND VGND VPWR VPWR _2980_ sky130_fd_sc_hd__clkbuf_1
X_4296_ _1762_ VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__clkbuf_1
X_3247_ _0795_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3178_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_83_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_1_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_37_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6937_ clknet_leaf_82_clk _0649_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cache_valid
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_91_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6868_ clknet_leaf_70_clk _0587_ net38 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_prediction\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5819_ tree_instances\[0\].u_tree.frame_id_out\[1\] tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[1\]
+ _0737_ VGND VGND VPWR VPWR _2848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_377 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6799_ clknet_leaf_42_clk _0521_ net33 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_208 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_463 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_321 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_68 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_105_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4150_ _1621_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6787__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4081_ _1555_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_37_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_102_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4983_ _1824_ _2229_ _2230_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__a21oi_1
XTAP_TAPCELL_ROW_34_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6722_ clknet_leaf_47_clk _0470_ net34 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_300 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_62_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3934_ _1413_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__clkbuf_1
X_6653_ clknet_leaf_32_clk _0017_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3865_ _1349_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6023__S _0799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5604_ _2576_ tree_instances\[8\].u_tree.frame_id_out\[0\] tree_instances\[8\].u_tree.frame_id_out\[2\]
+ _2619_ VGND VGND VPWR VPWR _2654_ sky130_fd_sc_hd__o22a_1
X_3796_ _1283_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__clkbuf_1
X_6584_ clknet_leaf_48_clk _0353_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5535_ _2590_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5466_ _2544_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4417_ _1850_ VGND VGND VPWR VPWR _1851_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_10_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_6_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5397_ _1136_ _2496_ _0006_ tree_instances\[10\].u_tree.pipeline_valid\[0\] VGND
+ VGND VPWR VPWR _0454_ sky130_fd_sc_hd__o2bb2a_1
X_4348_ _1803_ tree_instances\[5\].u_tree.pipeline_valid\[0\] tree_instances\[5\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__or3b_2
XFILLER_0_94_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4279_ _1746_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__clkbuf_1
X_6018_ tree_instances\[3\].u_tree.tree_state\[2\] tree_instances\[3\].u_tree.tree_state\[1\]
+ _2967_ VGND VGND VPWR VPWR _2971_ sky130_fd_sc_hd__or3_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_68_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__4388__S _0040_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6880__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_rst_buf_A rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_263 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_296 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_642 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_547 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3650_ tree_instances\[10\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1159_ sky130_fd_sc_hd__clkbuf_1
X_3581_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[2\] tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[3\]
+ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_11_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_2_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5320_ _1568_ _2414_ VGND VGND VPWR VPWR _2433_ sky130_fd_sc_hd__and2_1
X_5251_ _2396_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_458 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4202_ _1667_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5182_ _1355_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[3\] _2353_
+ _2354_ _2355_ VGND VGND VPWR VPWR _2356_ sky130_fd_sc_hd__o221a_1
XPHY_EDGE_ROW_79_Left_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4133_ _1589_ VGND VGND VPWR VPWR _1608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4064_ _1539_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6550__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xwire23 net9 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
XFILLER_0_64_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire12 _2689_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_19_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6705_ clknet_leaf_45_clk _0453_ net34 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_631 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4966_ tree_instances\[13\].u_tree.tree_state\[1\] _0967_ _1823_ VGND VGND VPWR VPWR
+ _2221_ sky130_fd_sc_hd__or3_1
XFILLER_0_61_303 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3917_ _1396_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__clkbuf_1
X_4897_ _1654_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[2\] _2169_
+ _2175_ _2176_ VGND VGND VPWR VPWR _2177_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_34_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6636_ clknet_leaf_32_clk _0395_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.current_node_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3848_ _1324_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__clkbuf_1
X_3779_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6567_ clknet_leaf_68_clk _0336_ net35 VGND VGND VPWR VPWR tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5518_ net2 _1020_ _2577_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__a21o_1
X_6498_ clknet_leaf_1_clk _0281_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ sky130_fd_sc_hd__dfxtp_1
X_5449_ _1492_ _2534_ VGND VGND VPWR VPWR _2536_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_74_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6638__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_311 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_92_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5723__A1 _2576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5723__B2 _2714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_408 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6379__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6308__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_88_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4820_ _1284_ _2071_ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_16_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_44_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4751_ tree_instances\[11\].u_tree.tree_state\[2\] tree_instances\[11\].u_tree.tree_state\[1\]
+ _1816_ VGND VGND VPWR VPWR _2070_ sky130_fd_sc_hd__or3_1
XFILLER_0_90_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_506 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3702_ _1202_ _1203_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__or2_1
XFILLER_0_83_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_54 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4682_ tree_instances\[10\].u_tree.read_enable VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__inv_2
X_3633_ _1142_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_99_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6421_ clknet_leaf_79_clk _0218_ VGND VGND VPWR VPWR tree_instances\[8\].u_tree.u_tree_weight_rom.gen_tree_8.u_tree_rom.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3564_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1083_ sky130_fd_sc_hd__clkbuf_1
X_6352_ clknet_leaf_20_clk _0159_ net25 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5303_ _2423_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__clkbuf_1
X_3495_ _1020_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6283_ _3141_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_110_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6731__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5234_ tree_instances\[17\].u_tree.frame_id_out\[4\] tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[4\]
+ tree_instances\[17\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_299 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5165_ _2338_ VGND VGND VPWR VPWR _2339_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4116_ _1590_ VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__clkbuf_1
X_5096_ tree_instances\[16\].u_tree.pipeline_prediction\[0\]\[0\] _2291_ _2293_ VGND
+ VGND VPWR VPWR _2294_ sky130_fd_sc_hd__mux2_1
X_4047_ _1523_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_203 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_78_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_439 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5998_ _2958_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_620 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4949_ _1718_ _2132_ VGND VGND VPWR VPWR _2211_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6619_ clknet_leaf_19_clk _0044_ net25 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_22_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6819__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5705__B2 _2598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6472__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6401__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_41_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_564 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_103_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3280_ _0822_ _0826_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__or2_1
X_6970_ clknet_leaf_81_clk _0676_ VGND VGND VPWR VPWR tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_5921_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[9\] _2900_ VGND VGND
+ VPWR VPWR _2911_ sky130_fd_sc_hd__and2_1
X_5852_ _1522_ _2426_ VGND VGND VPWR VPWR _2866_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5783_ complete_votes\[2\] VGND VGND VPWR VPWR _2826_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4803_ _1698_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[3\] VGND
+ VGND VPWR VPWR _2106_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_569 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4734_ _2061_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6983__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4665_ _2017_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3616_ tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1130_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6912__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4596_ _1972_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4340__A _1803_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6404_ clknet_leaf_91_clk _0206_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3547_ _1051_ _1058_ _1067_ tree_instances\[15\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0058_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6335_ clknet_leaf_93_clk _0143_ net27 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3478_ _1004_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__clkbuf_1
X_6266_ tree_instances\[5\].u_tree.current_node_data\[107\] tree_instances\[5\].u_tree.node_data\[107\]
+ _3132_ VGND VGND VPWR VPWR _3133_ sky130_fd_sc_hd__mux2_1
X_6197_ _3079_ _3034_ VGND VGND VPWR VPWR _3094_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_71_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5217_ _2379_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4674__A1 _1830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5148_ _0735_ _2322_ _0014_ tree_instances\[14\].u_tree.pipeline_valid\[0\] VGND
+ VGND VPWR VPWR _0378_ sky130_fd_sc_hd__o2bb2a_1
X_5079_ _2283_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_55_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6653__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_648 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_load_slew32_A tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_85_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_612 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6394__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_96_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4450_ _1877_ _1851_ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__and2_1
XFILLER_0_80_272 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4381_ _1825_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__inv_2
XANTENNA__6323__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3401_ _0935_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3332_ _0869_ _0873_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__or2_1
X_6120_ _3041_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6051_ _1247_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[6\] _2993_
+ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR VPWR _2994_
+ sky130_fd_sc_hd__a22o_1
X_3263_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _0810_ sky130_fd_sc_hd__clkbuf_1
X_3194_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__clkbuf_1
X_5002_ tree_instances\[13\].u_tree.read_enable VGND VGND VPWR VPWR _2240_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6953_ clknet_leaf_67_clk _0665_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[5\].u_tree.frame_id_out\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4335__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6884_ clknet_leaf_12_clk _0603_ net30 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_24_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5904_ _2902_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_5835_ tree_instances\[1\].u_tree.pipeline_prediction\[0\]\[0\] _2854_ _2857_ VGND
+ VGND VPWR VPWR _2858_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_52_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5766_ _2619_ tree_instances\[7\].u_tree.frame_id_out\[2\] tree_instances\[7\].u_tree.frame_id_out\[3\]
+ _2606_ VGND VGND VPWR VPWR _2811_ sky130_fd_sc_hd__a22o_1
X_5697_ _2603_ tree_instances\[17\].u_tree.frame_id_out\[1\] tree_instances\[17\].u_tree.frame_id_out\[3\]
+ _2659_ _2741_ VGND VGND VPWR VPWR _2742_ sky130_fd_sc_hd__a221oi_1
X_4717_ _2027_ tree_instances\[10\].u_tree.node_data\[12\] _2051_ tree_instances\[10\].u_tree.u_tree_weight_rom.gen_tree_10.u_tree_rom.node_data\[12\]
+ VGND VGND VPWR VPWR _2052_ sky130_fd_sc_hd__a22o_1
X_4648_ _1598_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[3\] tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ _1581_ VGND VGND VPWR VPWR _2006_ sky130_fd_sc_hd__a2bb2o_1
XPHY_EDGE_ROW_15_Left_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4579_ _1799_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[5\] _1956_
+ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_93 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6318_ clknet_leaf_15_clk _0127_ net28 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
X_6249_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[7\] _2475_ _3116_
+ VGND VGND VPWR VPWR _3124_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_24_Left_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_4_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_80_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6834__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_401 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_33_Left_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_91_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_18 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_42_Left_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3950_ _1401_ _0771_ _1426_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__and3_1
XFILLER_0_85_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3881_ _1222_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6575__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_51_Left_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5620_ _2602_ tree_instances\[12\].u_tree.frame_id_out\[1\] _2668_ _2582_ _2669_
+ VGND VGND VPWR VPWR _2670_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_100_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_209 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6504__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5551_ _2598_ tree_instances\[20\].u_tree.frame_id_out\[0\] tree_instances\[20\].u_tree.frame_id_out\[2\]
+ _2600_ VGND VGND VPWR VPWR _2601_ sky130_fd_sc_hd__o2bb2a_1
X_4502_ _1310_ _1840_ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_294 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_369 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5482_ _2554_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4433_ _1863_ _1851_ VGND VGND VPWR VPWR _1864_ sky130_fd_sc_hd__and2_1
XANTENNA__5714__A _2622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4364_ _1112_ tree_instances\[11\].u_tree.pipeline_valid\[0\] tree_instances\[11\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__or3b_2
X_6103_ _3031_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_60_Left_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_597 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4295_ _1037_ VGND VGND VPWR VPWR _1762_ sky130_fd_sc_hd__clkbuf_1
X_3315_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0858_ sky130_fd_sc_hd__clkbuf_1
X_6034_ _2872_ _2517_ VGND VGND VPWR VPWR _2979_ sky130_fd_sc_hd__nor2_1
X_3246_ _0792_ _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__nor2_1
X_3177_ _0731_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__buf_4
XFILLER_0_83_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_1_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6936_ clknet_leaf_94_clk _0648_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_prediction\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_180 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_76_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6867_ clknet_leaf_17_clk _0586_ net28 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6798_ clknet_leaf_41_clk _0520_ net33 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_5818_ _2847_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5749_ tree_instances\[11\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2794_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5624__A _2610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_9_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_345 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4080_ _1554_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6756__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4982_ _1114_ _1824_ VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__nor2_1
X_6721_ clknet_leaf_34_clk _0469_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_62_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_98 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3933_ _0764_ VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6652_ clknet_leaf_35_clk _0059_ net33 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_73_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3864_ _1195_ _1337_ _1348_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5603_ tree_instances\[13\].u_tree.prediction_out _2645_ _2652_ tree_instances\[1\].u_tree.prediction_out
+ VGND VGND VPWR VPWR _2653_ sky130_fd_sc_hd__a22o_1
X_6583_ clknet_leaf_48_clk _0352_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3795_ _1203_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5534_ _2589_ net6 _1020_ VGND VGND VPWR VPWR _2590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5465_ tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[1\] _2246_ _0028_ VGND
+ VGND VPWR VPWR _2544_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4416_ tree_instances\[6\].u_tree.tree_state\[1\] tree_instances\[6\].u_tree.tree_state\[2\]
+ _1811_ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__or3_1
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_6_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_372 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5396_ tree_instances\[10\].u_tree.tree_state\[0\] tree_instances\[10\].u_tree.pipeline_valid\[0\]
+ VGND VGND VPWR VPWR _2496_ sky130_fd_sc_hd__nand2_1
X_4347_ _1807_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__inv_2
XFILLER_0_94_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5275__A1 _2246_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4278_ _1736_ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3229_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__clkbuf_1
X_6017_ tree_instances\[3\].u_tree.tree_state\[0\] _0851_ tree_instances\[3\].u_tree.tree_state\[1\]
+ VGND VGND VPWR VPWR _2970_ sky130_fd_sc_hd__o21ba_1
XTAP_TAPCELL_ROW_68_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6919_ clknet_leaf_24_clk _0632_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.frame_id_out\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_472 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_24_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_79_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_141 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_82_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_13 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5529__A _2585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_97_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_559 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3580_ tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[0\] tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[1\]
+ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_3_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_11_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5250_ _1385_ _2313_ VGND VGND VPWR VPWR _2396_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4201_ _1672_ VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__clkbuf_1
X_5181_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[5\] tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ VGND VGND VPWR VPWR _2355_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4701__B1 _0010_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4132_ _1605_ VGND VGND VPWR VPWR _1607_ sky130_fd_sc_hd__clkbuf_1
X_4063_ _1529_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xwire13 net14 VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6590__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_19_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4965_ tree_instances\[13\].u_tree.tree_state\[1\] _2166_ VGND VGND VPWR VPWR _2220_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_120 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3916_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1396_ sky130_fd_sc_hd__clkbuf_1
X_6704_ clknet_leaf_83_clk _0452_ net31 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4896_ _0962_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[4\] VGND
+ VGND VPWR VPWR _2176_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6635_ clknet_leaf_62_clk _0394_ net37 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3847_ _1192_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_389 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3778_ _1267_ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6566_ clknet_leaf_21_clk _0082_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5517_ _2576_ _1019_ VGND VGND VPWR VPWR _2577_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_14_275 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6497_ clknet_leaf_1_clk _0280_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[6\]
+ sky130_fd_sc_hd__dfxtp_1
X_5448_ _2535_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_74_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5379_ _2480_ VGND VGND VPWR VPWR _2481_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6678__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6607__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_29_Right_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_7_Left_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_EDGE_ROW_38_Right_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_47_Right_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_88_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6348__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_312 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_44_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_56_Right_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4750_ _2069_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__clkbuf_1
X_3701_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_518 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4681_ _2025_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__clkbuf_1
X_3632_ _1141_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND
+ VPWR VPWR _1142_ sky130_fd_sc_hd__or2_1
XTAP_TAPCELL_ROW_99_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6420_ clknet_leaf_94_clk _0217_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5706__B _2578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6351_ clknet_leaf_20_clk _0158_ net25 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_3563_ tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1082_ sky130_fd_sc_hd__clkbuf_1
X_5302_ tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[2\] _2125_ _0024_ VGND
+ VGND VPWR VPWR _2423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3494_ _1019_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6282_ _2481_ _3102_ VGND VGND VPWR VPWR _3141_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_110_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_65_Right_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5233_ _2387_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__clkbuf_1
X_5164_ _2337_ VGND VGND VPWR VPWR _2338_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5722__A _2714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4115_ _1583_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6771__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5095_ tree_instances\[16\].u_tree.tree_state\[0\] _1022_ _0017_ _2292_ VGND VGND
+ VPWR VPWR _2293_ sky130_fd_sc_hd__a211oi_1
X_4046_ _1518_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_EDGE_ROW_74_Right_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5997_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[5\] _1424_ _2899_
+ VGND VGND VPWR VPWR _2958_ sky130_fd_sc_hd__mux2_1
X_4948_ _2210_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_602 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4879_ _2154_ VGND VGND VPWR VPWR _2160_ sky130_fd_sc_hd__clkbuf_1
X_6618_ clknet_leaf_20_clk _0043_ net24 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5616__B _2585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6549_ clknet_leaf_42_clk _0323_ net36 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_83_Right_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5469__A1 _2249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6859__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6441__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_234 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_92_Right_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_418 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_553 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_65_473 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_145 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5632__A1 _2606_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5920_ _2910_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5851_ _2865_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_100_Right_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5782_ _2824_ _2825_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__nor2_1
X_4802_ _1702_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND
+ VGND VPWR VPWR _2105_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4733_ _1610_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[6\] _2010_
+ VGND VGND VPWR VPWR _2061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4664_ _1639_ _2012_ VGND VGND VPWR VPWR _2017_ sky130_fd_sc_hd__and2_1
XANTENNA__5699__A1 _2659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6403_ clknet_leaf_9_clk _0205_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3615_ tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1129_ sky130_fd_sc_hd__clkbuf_1
X_4595_ tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[3\] _1835_ _0044_ VGND
+ VGND VPWR VPWR _1972_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3546_ _1064_ _1066_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__nor2_1
XFILLER_0_3_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6334_ clknet_leaf_90_clk _0142_ net27 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6952__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6265_ _0933_ VGND VGND VPWR VPWR _3132_ sky130_fd_sc_hd__clkbuf_1
X_3477_ _1002_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__or2_1
X_5216_ tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[1\] _2246_ _0020_ VGND
+ VGND VPWR VPWR _2379_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6196_ _3093_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5147_ tree_instances\[14\].u_tree.pipeline_valid\[0\] tree_instances\[14\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _2322_ sky130_fd_sc_hd__nand2_1
X_5078_ _1542_ _2255_ VGND VGND VPWR VPWR _2283_ sky130_fd_sc_hd__and2_1
X_4029_ _0884_ VGND VGND VPWR VPWR _1506_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_55_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_27_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_66_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5627__A _2582_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_97_Left_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6693__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6622__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5862__A1 tree_instances\[0\].u_tree.frame_id_in\[4\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_89_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_85_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5614__A1 _2600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_624 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_432 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5537__A _1827_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4380_ _1112_ tree_instances\[19\].u_tree.pipeline_valid\[0\] tree_instances\[19\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__or3b_1
X_3400_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[0\] tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[1\]
+ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__or2_1
X_3331_ _0871_ _0872_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6050_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[7\] VGND VGND VPWR
+ VPWR _2993_ sky130_fd_sc_hd__inv_2
X_3262_ _0803_ _0806_ _0807_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__o211a_1
X_3193_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _0746_ sky130_fd_sc_hd__buf_1
X_5001_ _2239_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6525__SET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5605__A1 _2575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6952_ clknet_leaf_83_clk _0664_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.read_enable
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5903_ _2147_ _2901_ VGND VGND VPWR VPWR _2902_ sky130_fd_sc_hd__and2_1
X_6883_ clknet_leaf_71_clk _0602_ net38 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.read_enable
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5834_ _1821_ net17 _2855_ _2856_ VGND VGND VPWR VPWR _2857_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_52_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_24_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_309 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5765_ _2804_ _2806_ _2809_ VGND VGND VPWR VPWR _2810_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_123 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5696_ _2582_ tree_instances\[17\].u_tree.frame_id_out\[2\] VGND VGND VPWR VPWR _2741_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_156 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4716_ _2050_ VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4647_ _1994_ _2002_ _2003_ _2004_ VGND VGND VPWR VPWR _2005_ sky130_fd_sc_hd__or4bb_1
X_6317_ clknet_leaf_30_clk _0126_ net28 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_4578_ _1962_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3529_ _1034_ _1038_ _1045_ _1050_ tree_instances\[8\].u_tree.tree_state\[1\] VGND
+ VGND VPWR VPWR _0084_ sky130_fd_sc_hd__a41o_1
XFILLER_0_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6248_ _3123_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__clkbuf_1
X_6179_ _3085_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_4_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_240 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6803__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_91_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_35 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3880_ _0918_ _0924_ _0930_ _1359_ _1363_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a32o_1
Xclkbuf_leaf_70_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA__6012__A1 tree_instances\[0\].u_tree.frame_id_in\[4\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_100_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5550_ _2599_ VGND VGND VPWR VPWR _2600_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_100_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4501_ _1920_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5481_ tree_instances\[20\].u_tree.frame_id_out\[0\] tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _1197_ VGND VGND VPWR VPWR _2554_ sky130_fd_sc_hd__mux2_1
X_4432_ _1862_ VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6544__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_521 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4363_ _1815_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__buf_2
X_6102_ tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[4\] tree_instances\[0\].u_tree.frame_id_in\[4\]
+ _0034_ VGND VGND VPWR VPWR _3031_ sky130_fd_sc_hd__mux2_1
X_4294_ _1761_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_3314_ _0856_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__clkbuf_1
X_3245_ _0793_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__clkbuf_1
X_6033_ _0799_ _0800_ _2967_ tree_instances\[3\].u_tree.ready_for_next VGND VGND VPWR
+ VPWR _0609_ sky130_fd_sc_hd__a22o_1
X_3176_ _0730_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__buf_4
XANTENNA__4346__A _1803_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_1_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6935_ clknet_leaf_31_clk _0647_ net33 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_65_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_4
X_6866_ clknet_leaf_40_clk _0100_ net30 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5817_ tree_instances\[0\].u_tree.frame_id_out\[0\] tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[0\]
+ _0737_ VGND VGND VPWR VPWR _2847_ sky130_fd_sc_hd__mux2_1
X_6797_ clknet_leaf_98_clk _0052_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_107_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_106_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5748_ _2576_ tree_instances\[11\].u_tree.frame_id_out\[0\] tree_instances\[11\].u_tree.frame_id_out\[2\]
+ _2619_ _2792_ VGND VGND VPWR VPWR _2793_ sky130_fd_sc_hd__o221a_1
XFILLER_0_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5679_ _2586_ tree_instances\[4\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2724_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_3_5__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_392 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_32_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5640__A _2614_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__7002__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_52_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_593 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_93_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput2 net2 VGND VGND VPWR VPWR frame_id_out[0] sky130_fd_sc_hd__buf_8
XFILLER_0_77_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4981_ _1822_ _1114_ tree_instances\[13\].u_tree.ready_for_next VGND VGND VPWR VPWR
+ _2229_ sky130_fd_sc_hd__a21oi_1
X_6720_ clknet_leaf_48_clk _0468_ net34 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_102_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_62_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3932_ _1177_ _1394_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_34_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_184 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6651_ clknet_leaf_66_clk _0095_ net36 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4613__B _1937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6796__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3863_ _1324_ _1340_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__nor2_1
X_6582_ clknet_leaf_48_clk _0351_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6725__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5602_ _2646_ _2648_ _2651_ VGND VGND VPWR VPWR _2652_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_613 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_5_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3794_ _1282_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__clkbuf_1
X_5533_ _2588_ VGND VGND VPWR VPWR _2589_ sky130_fd_sc_hd__buf_4
XFILLER_0_6_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5464_ _2543_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4415_ _1848_ VGND VGND VPWR VPWR _1849_ sky130_fd_sc_hd__clkbuf_1
X_5395_ _0737_ _2495_ _0004_ tree_instances\[0\].u_tree.pipeline_valid\[0\] VGND VGND
+ VPWR VPWR _0453_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4346_ _1803_ tree_instances\[4\].u_tree.pipeline_valid\[0\] tree_instances\[4\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__or3b_2
XTAP_TAPCELL_ROW_6_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4277_ _1744_ VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__clkbuf_1
X_3228_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[8\] tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[7\]
+ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__nor2_1
X_6016_ _2968_ VGND VGND VPWR VPWR _2969_ sky130_fd_sc_hd__clkbuf_1
X_3159_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _0715_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_4
X_6918_ clknet_leaf_23_clk _0631_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.frame_id_out\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6849_ clknet_leaf_40_clk _0569_ net36 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6466__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_221 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_153 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_25_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_140 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_max_cap29_A net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_36_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4200_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1672_ sky130_fd_sc_hd__clkbuf_1
X_5180_ _1217_ tree_instances\[16\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND
+ VGND VPWR VPWR _2354_ sky130_fd_sc_hd__and2_1
XFILLER_0_48_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4131_ _1599_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__clkbuf_1
X_4062_ _1532_ VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire14 net16 VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
XANTENNA__6977__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_19_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_47_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_16_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4964_ _2218_ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__clkbuf_1
X_6703_ clknet_leaf_7_clk _0451_ net25 VGND VGND VPWR VPWR state\[1\] sky130_fd_sc_hd__dfrtp_1
X_3915_ _1173_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_132 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4895_ _1656_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[0\] VGND
+ VGND VPWR VPWR _2175_ sky130_fd_sc_hd__nor2_1
X_6634_ clknet_leaf_62_clk _0393_ net35 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3846_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1331_ sky130_fd_sc_hd__clkbuf_1
X_3777_ _1141_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6565_ clknet_leaf_21_clk _0040_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6496_ clknet_leaf_102_clk _0279_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[5\]
+ sky130_fd_sc_hd__dfxtp_1
X_5516_ _2575_ VGND VGND VPWR VPWR _2576_ sky130_fd_sc_hd__buf_4
X_5447_ _1496_ _2534_ VGND VGND VPWR VPWR _2535_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5378_ _0940_ VGND VGND VPWR VPWR _2480_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_74_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4329_ _1775_ _1782_ VGND VGND VPWR VPWR _1796_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6647__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_121 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_165 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_16_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6388__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_44_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6317__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3700_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__clkbuf_1
X_4680_ tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[4\] _1837_ _0006_ VGND
+ VGND VPWR VPWR _2025_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3631_ tree_instances\[11\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1141_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_124 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_70_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3562_ _1072_ _1074_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_99_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6350_ clknet_leaf_20_clk _0157_ net25 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5301_ _2422_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_574 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3493_ state\[0\] _1018_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__or2_1
X_6281_ _3140_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_110_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5232_ tree_instances\[17\].u_tree.frame_id_out\[3\] tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[3\]
+ _0909_ VGND VGND VPWR VPWR _2387_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_268 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_5_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_4
X_5163_ _0792_ VGND VGND VPWR VPWR _2337_ sky130_fd_sc_hd__clkbuf_1
X_4114_ _1588_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__clkbuf_1
X_5094_ tree_instances\[16\].u_tree.tree_state\[1\] tree_instances\[16\].u_tree.tree_state\[2\]
+ tree_instances\[16\].u_tree.tree_state\[0\] VGND VGND VPWR VPWR _2292_ sky130_fd_sc_hd__nor3_1
X_4045_ _1521_ VGND VGND VPWR VPWR _1522_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4354__A _1803_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6740__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5996_ _2957_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4947_ _1726_ _2133_ VGND VGND VPWR VPWR _2210_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4878_ _2150_ VGND VGND VPWR VPWR _2159_ sky130_fd_sc_hd__clkbuf_1
X_3829_ _0951_ tree_instances\[11\].u_tree.prediction_valid VGND VGND VPWR VPWR _0089_
+ sky130_fd_sc_hd__nor2_1
X_6617_ clknet_leaf_19_clk _0085_ net25 VGND VGND VPWR VPWR tree_instances\[9\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6548_ clknet_leaf_45_clk _0322_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_76_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_81_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6479_ clknet_leaf_10_clk _0267_ net25 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_96_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6828__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6481__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_97_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6700__SET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6410__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_622 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_34_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_41_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_565 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_49_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_21_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_405 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_49_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6569__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap1 net42 VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
X_5850_ _1510_ _2427_ VGND VGND VPWR VPWR _2865_ sky130_fd_sc_hd__and2_1
XFILLER_0_68_290 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5781_ _2729_ _2820_ _1018_ complete_votes\[1\] complete_votes\[0\] VGND VGND VPWR
+ VPWR _2825_ sky130_fd_sc_hd__o2111a_1
X_4801_ _1691_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[5\] VGND
+ VGND VPWR VPWR _2104_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_69 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_83_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4732_ _2060_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__clkbuf_1
X_4663_ _2016_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3614_ _1125_ _1127_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__nor2_1
XANTENNA__4621__B _1937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6402_ clknet_leaf_91_clk _0204_ net27 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4594_ _1971_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_1
X_3545_ _1065_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6333_ clknet_leaf_91_clk _0141_ net27 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_6264_ _3131_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__clkbuf_1
X_3476_ tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1003_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5215_ _2378_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__clkbuf_1
X_6195_ _2563_ _3034_ VGND VGND VPWR VPWR _3093_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_71_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3253__A _0799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5146_ _1023_ _2321_ _1809_ tree_instances\[16\].u_tree.ready_for_next VGND VGND
+ VPWR VPWR _0377_ sky130_fd_sc_hd__a22o_1
XANTENNA__6992__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5077_ _2282_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6921__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4028_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1505_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5979_ _1335_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[6\] _2944_
+ _2945_ VGND VGND VPWR VPWR _2946_ sky130_fd_sc_hd__o211a_1
XTAP_TAPCELL_ROW_82_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_282 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_62_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_514 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_57_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_395 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_96_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_505 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3330_ tree_instances\[1\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _0872_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5302__A1 _2125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3261_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[9\] VGND VGND VPWR
+ VPWR _0808_ sky130_fd_sc_hd__inv_2
X_5000_ _1673_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[7\] _2189_
+ VGND VGND VPWR VPWR _2239_ sky130_fd_sc_hd__mux2_1
X_3192_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _0745_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6332__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_43 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6951_ clknet_leaf_90_clk _0663_ net31 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_105_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5902_ _2900_ VGND VGND VPWR VPWR _2901_ sky130_fd_sc_hd__dlymetal6s2s_1
X_6882_ clknet_leaf_89_clk _0601_ net30 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5833_ tree_instances\[1\].u_tree.tree_state\[1\] tree_instances\[1\].u_tree.tree_state\[0\]
+ tree_instances\[1\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _2856_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5764_ _2619_ tree_instances\[6\].u_tree.frame_id_out\[2\] _2807_ _2589_ _2808_ VGND
+ VGND VPWR VPWR _2809_ sky130_fd_sc_hd__o221a_1
XFILLER_0_56_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5695_ _2576_ tree_instances\[17\].u_tree.frame_id_out\[0\] tree_instances\[17\].u_tree.frame_id_out\[1\]
+ _2713_ VGND VGND VPWR VPWR _2740_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4715_ _2049_ VGND VGND VPWR VPWR _2050_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4646_ _1599_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[3\] VGND
+ VGND VPWR VPWR _2004_ sky130_fd_sc_hd__nand2_1
XFILLER_0_16_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4577_ _1800_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[4\] _1956_
+ VGND VGND VPWR VPWR _1962_ sky130_fd_sc_hd__mux2_1
XANTENNA_wire1_A clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6316_ clknet_leaf_30_clk _0125_ net28 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3528_ _1048_ _1049_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__nor2_1
X_3459_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[8\] VGND VGND VPWR
+ VPWR _0989_ sky130_fd_sc_hd__clkbuf_1
X_6247_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[6\] _2474_ _3116_
+ VGND VGND VPWR VPWR _3123_ sky130_fd_sc_hd__mux2_1
X_6178_ tree_instances\[5\].u_tree.pipeline_prediction\[0\]\[0\] _3082_ _3084_ VGND
+ VGND VPWR VPWR _3085_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5129_ tree_instances\[16\].u_tree.tree_state\[1\] _2292_ VGND VGND VPWR VPWR _2312_
+ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_4_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_436 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_31_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6843__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_138 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5548__A _2575_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5771__A1 _2713_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_241 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_26_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4500_ _1304_ _1840_ VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5480_ _2502_ _2551_ _2553_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__a21bo_1
X_4431_ _1861_ VGND VGND VPWR VPWR _1862_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_1 tree_instances\[13\].u_tree.prediction_out VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_22_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4362_ tree_instances\[15\].u_tree.pipeline_valid\[0\] tree_instances\[15\].u_tree.tree_state\[0\]
+ net1 VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__and3b_1
XANTENNA__6584__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4293_ tree_instances\[6\].u_tree.prediction_valid _0932_ VGND VGND VPWR VPWR _1761_
+ sky130_fd_sc_hd__and2b_1
X_6101_ _3030_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__clkbuf_1
X_3313_ _0855_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND
+ VPWR VPWR _0856_ sky130_fd_sc_hd__or2_1
X_3244_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _0793_ sky130_fd_sc_hd__buf_1
XANTENNA__6513__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6032_ _2978_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__clkbuf_1
X_3175_ net1 VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_1_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6934_ clknet_leaf_74_clk _0646_ VGND VGND VPWR VPWR tree_instances\[20\].u_tree.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XTAP_TAPCELL_ROW_37_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_65_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6865_ clknet_leaf_67_clk _0585_ net36 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_49_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5816_ _2846_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_76_388 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_539 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_8_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6796_ clknet_leaf_98_clk _0010_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5747_ _2586_ tree_instances\[11\].u_tree.frame_id_out\[3\] VGND VGND VPWR VPWR _2792_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_230 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5678_ _2589_ tree_instances\[4\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2723_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4629_ tree_instances\[19\].u_tree.tree_state\[0\] _1251_ VGND VGND VPWR VPWR _1989_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_9_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5640__B _2636_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_620 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_93_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput3 net3 VGND VGND VPWR VPWR frame_id_out[1] sky130_fd_sc_hd__buf_8
XFILLER_0_37_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4980_ _2228_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_102_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3931_ _1404_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_34_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_196 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6650_ clknet_leaf_57_clk _0409_ net37 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
X_3862_ _1321_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6581_ clknet_leaf_48_clk _0350_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_5601_ _2575_ tree_instances\[1\].u_tree.frame_id_out\[0\] tree_instances\[1\].u_tree.prediction_valid
+ _2649_ _2650_ VGND VGND VPWR VPWR _2651_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_6_625 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_39_591 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3793_ _1201_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_550 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5532_ current_voting_frame\[4\] VGND VGND VPWR VPWR _2588_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6765__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5463_ tree_instances\[20\].u_tree.pipeline_frame_id\[0\]\[0\] _2122_ _0028_ VGND
+ VGND VPWR VPWR _2543_ sky130_fd_sc_hd__mux2_1
X_4414_ _1847_ VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__clkbuf_1
X_5394_ tree_instances\[0\].u_tree.tree_state\[0\] _0736_ VGND VGND VPWR VPWR _2495_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4345_ _1806_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_6_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5741__A _2627_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4276_ _1730_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_85 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3227_ _0775_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__clkbuf_1
X_6015_ tree_instances\[3\].u_tree.read_enable VGND VGND VPWR VPWR _2968_ sky130_fd_sc_hd__inv_2
X_3158_ tree_instances\[4\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _0714_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_68_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6917_ clknet_leaf_17_clk _0630_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6848_ clknet_leaf_40_clk _0568_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6779_ clknet_leaf_7_clk _0513_ net25 VGND VGND VPWR VPWR complete_votes\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_79_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_233 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5635__B _2579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6435__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_347 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_82_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_11_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_11_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_39_Left_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6650__SET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4130_ _1597_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5561__A _2610_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4061_ _1530_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_48_Left_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_19_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4963_ tree_instances\[13\].u_tree.read_enable VGND VGND VPWR VPWR _2218_ sky130_fd_sc_hd__inv_2
XTAP_TAPCELL_ROW_47_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_65 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3914_ _1393_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__clkbuf_1
X_6702_ clknet_leaf_7_clk _0450_ net25 VGND VGND VPWR VPWR state\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5717__A1 _2619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6633_ clknet_leaf_64_clk _0392_ net35 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4894_ _2172_ _2173_ VGND VGND VPWR VPWR _2174_ sky130_fd_sc_hd__nand2_1
XANTENNA__6946__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5717__B2 _2586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3845_ _1187_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3776_ _1154_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__clkbuf_1
X_6564_ clknet_leaf_21_clk _0039_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6495_ clknet_leaf_101_clk _0278_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_6_488 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5515_ current_voting_frame\[0\] VGND VGND VPWR VPWR _2575_ sky130_fd_sc_hd__inv_2
X_5446_ _2533_ VGND VGND VPWR VPWR _2534_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5377_ _1240_ _2471_ VGND VGND VPWR VPWR _2479_ sky130_fd_sc_hd__nand2_1
XTAP_TAPCELL_ROW_74_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4328_ _1794_ VGND VGND VPWR VPWR _1795_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_input1_A feature_valid VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4259_ tree_instances\[5\].u_tree.prediction_valid _0903_ VGND VGND VPWR VPWR _1728_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_417 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_84_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6687__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_177 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_52_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_269 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_8_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6786__SET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3630_ tree_instances\[11\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3561_ _1072_ _1074_ _1076_ _1079_ _1080_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__o41a_1
X_5300_ tree_instances\[19\].u_tree.pipeline_frame_id\[0\]\[1\] _2246_ _0024_ VGND
+ VGND VPWR VPWR _2422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3492_ state\[1\] VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__inv_2
X_6280_ _2486_ _3102_ VGND VGND VPWR VPWR _3140_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_110_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5231_ _2386_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__clkbuf_1
X_5162_ _2335_ VGND VGND VPWR VPWR _2336_ sky130_fd_sc_hd__clkbuf_1
X_5093_ tree_instances\[16\].u_tree.tree_state\[1\] tree_instances\[16\].u_tree.current_node_data\[12\]
+ tree_instances\[16\].u_tree.node_data\[12\] _2290_ VGND VGND VPWR VPWR _2291_ sky130_fd_sc_hd__a22o_1
XANTENNA__4619__B _1937_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4113_ _1587_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4044_ _1228_ VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5995_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[4\] _1421_ _2899_
+ VGND VGND VPWR VPWR _2957_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4946_ _2209_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6780__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4877_ _2140_ VGND VGND VPWR VPWR _2158_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6616_ clknet_leaf_93_clk _0379_ VGND VGND VPWR VPWR tree_instances\[10\].u_tree.u_tree_weight_rom.gen_tree_10.u_tree_rom.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XANTENNA__4370__A _1112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_380 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3828_ _1315_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6547_ clknet_leaf_3_clk _0321_ net26 VGND VGND VPWR VPWR tree_instances\[13\].u_tree.current_node_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3759_ tree_instances\[19\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_76_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_501 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_400 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6478_ clknet_leaf_9_clk _0266_ net27 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5429_ _1497_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[3\] _2519_
+ VGND VGND VPWR VPWR _2523_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_280 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_97_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_512 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5929__A1 _1834_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6868__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_41_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6450__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_21_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_36 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_49_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_29_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_61_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4800_ _2100_ _2101_ _2102_ VGND VGND VPWR VPWR _2103_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_67 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5780_ _2447_ _2707_ _2821_ _0000_ _2823_ VGND VGND VPWR VPWR _2824_ sky130_fd_sc_hd__o32a_1
X_4731_ _1614_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[5\] _2010_
+ VGND VGND VPWR VPWR _2060_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4662_ _1633_ _2012_ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3613_ _1126_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6401_ clknet_leaf_91_clk _0203_ net25 VGND VGND VPWR VPWR tree_instances\[10\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4593_ tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[2\] _1832_ _0044_ VGND
+ VGND VPWR VPWR _1971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3544_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[1\] tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[2\]
+ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__or2_1
X_6332_ clknet_leaf_90_clk _0140_ net31 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_6263_ tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[4\] tree_instances\[0\].u_tree.frame_id_in\[4\]
+ _0038_ VGND VGND VPWR VPWR _3131_ sky130_fd_sc_hd__mux2_1
X_3475_ tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _1002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5214_ tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[0\] _2122_ _0020_ VGND
+ VGND VPWR VPWR _2378_ sky130_fd_sc_hd__mux2_1
X_6194_ _3092_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5145_ tree_instances\[16\].u_tree.tree_state\[0\] _1022_ VGND VGND VPWR VPWR _2321_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5076_ _1546_ _2255_ VGND VGND VPWR VPWR _2282_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4027_ _1503_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4831__A1 _1830_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5978_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[0\] _2939_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[1\]
+ _1322_ tree_instances\[3\].u_tree.u_tree_weight_rom.cache_valid VGND VGND VPWR VPWR
+ _2945_ sky130_fd_sc_hd__o221a_1
XTAP_TAPCELL_ROW_82_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5599__B_N _2585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4929_ _2200_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_489 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_375 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_89_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_26_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6631__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_54_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_96_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_111_517 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_236 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3260_ tree_instances\[2\].u_tree.pipeline_current_node\[0\]\[8\] VGND VGND VPWR
+ VPWR _0807_ sky130_fd_sc_hd__inv_2
X_3191_ _0743_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND
+ VPWR VPWR _0744_ sky130_fd_sc_hd__or2_1
XFILLER_0_56_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6950_ clknet_leaf_87_clk _0662_ net30 VGND VGND VPWR VPWR tree_instances\[5\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6719__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_80_clk_A clknet_3_4__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5901_ tree_instances\[2\].u_tree.tree_state\[2\] tree_instances\[2\].u_tree.tree_state\[1\]
+ _1804_ VGND VGND VPWR VPWR _2900_ sky130_fd_sc_hd__or3_1
XTAP_TAPCELL_ROW_105_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6881_ clknet_leaf_13_clk _0600_ net29 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5832_ tree_instances\[1\].u_tree.tree_state\[0\] _1226_ VGND VGND VPWR VPWR _2855_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_548 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6372__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5763_ _2600_ tree_instances\[6\].u_tree.frame_id_out\[2\] tree_instances\[6\].u_tree.frame_id_out\[3\]
+ _2606_ VGND VGND VPWR VPWR _2808_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__6301__RESET_B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_336 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_56_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4714_ tree_instances\[10\].u_tree.read_enable _2008_ VGND VGND VPWR VPWR _2049_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_16_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5694_ tree_instances\[17\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2739_ sky130_fd_sc_hd__inv_2
XFILLER_0_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4645_ _1159_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[2\] VGND
+ VGND VPWR VPWR _2003_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4576_ _1961_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6315_ clknet_leaf_24_clk _0124_ net28 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_342 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3527_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1049_ sky130_fd_sc_hd__buf_1
XANTENNA_clkbuf_leaf_33_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3458_ _0976_ _0987_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__nor2_1
X_6246_ _3122_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__clkbuf_1
X_3389_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND VPWR
+ VPWR _0926_ sky130_fd_sc_hd__buf_1
XANTENNA_wire22_A net23 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6177_ tree_instances\[5\].u_tree.tree_state\[0\] _0902_ _0035_ _3083_ VGND VGND
+ VPWR VPWR _3084_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_99_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5128_ _2310_ VGND VGND VPWR VPWR _2311_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5057__A1 _2125_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_48_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_84_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5059_ tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[3\] _2249_ _0016_ VGND
+ VGND VPWR VPWR _2273_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_79_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_51_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_109_Right_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6883__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_load_slew30_A tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_11_Left_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_529 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5220__A1 _2249_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_100_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4430_ _1860_ VGND VGND VPWR VPWR _1861_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_20_Left_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6100_ tree_instances\[4\].u_tree.pipeline_frame_id\[0\]\[3\] _1834_ _0034_ VGND
+ VGND VPWR VPWR _3030_ sky130_fd_sc_hd__mux2_1
X_4361_ _1814_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_545 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4292_ _1734_ VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__clkbuf_1
X_3312_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _0855_ sky130_fd_sc_hd__clkbuf_1
X_3243_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _0792_ sky130_fd_sc_hd__buf_1
X_6031_ tree_instances\[3\].u_tree.prediction_out tree_instances\[3\].u_tree.pipeline_prediction\[0\]\[0\]
+ tree_instances\[3\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2978_ sky130_fd_sc_hd__mux2_1
X_3174_ _0709_ _0721_ _0728_ _0729_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__o31a_1
XFILLER_0_83_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6553__RESET_B net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_1_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6933_ clknet_leaf_36_clk _0645_ net33 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5739__A _2579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_65_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6864_ clknet_leaf_69_clk _0584_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_TAPCELL_ROW_37_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5815_ tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[4\] _2251_ _0004_ VGND
+ VGND VPWR VPWR _2846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6795_ clknet_leaf_99_clk _0009_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.tree_state\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5746_ _2576_ tree_instances\[11\].u_tree.frame_id_out\[0\] _2789_ _2790_ VGND VGND
+ VPWR VPWR _2791_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_57_592 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5677_ _2589_ tree_instances\[4\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2722_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_44_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4628_ _1025_ _1988_ _1814_ tree_instances\[9\].u_tree.ready_for_next VGND VGND VPWR
+ VPWR _0191_ sky130_fd_sc_hd__a22o_1
X_4559_ _1952_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_9_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6229_ _2310_ _2360_ VGND VGND VPWR VPWR _3112_ sky130_fd_sc_hd__nor2_1
XTAP_TAPCELL_ROW_90_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_632 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_93_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xoutput4 net4 VGND VGND VPWR VPWR frame_id_out[2] sky130_fd_sc_hd__buf_8
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3930_ _1409_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5559__A _2578_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_102_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_46_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3861_ _1345_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6580_ clknet_leaf_49_clk _0349_ net35 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_current_node\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3792_ _1277_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5600_ _2610_ tree_instances\[1\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2650_
+ sky130_fd_sc_hd__xnor2_1
X_5531_ _2587_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_562 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_201 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5462_ _2542_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4413_ _1846_ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__clkbuf_1
X_5393_ _1000_ _2494_ _0042_ tree_instances\[8\].u_tree.pipeline_valid\[0\] VGND VGND
+ VPWR VPWR _0452_ sky130_fd_sc_hd__o2bb2a_1
X_4344_ tree_instances\[3\].u_tree.pipeline_valid\[0\] tree_instances\[3\].u_tree.tree_state\[0\]
+ net1 VGND VGND VPWR VPWR _1806_ sky130_fd_sc_hd__and3b_1
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_6_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_492 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4275_ _1731_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__clkbuf_1
X_6014_ _0032_ VGND VGND VPWR VPWR _2967_ sky130_fd_sc_hd__inv_2
XANTENNA__6734__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5680__A1 _2576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3226_ tree_instances\[17\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_97 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3157_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5680__B2 _2714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_68_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6916_ clknet_leaf_17_clk _0629_ net28 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.frame_id_out\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6847_ clknet_leaf_89_clk _0567_ net30 VGND VGND VPWR VPWR tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6778_ clknet_leaf_6_clk _0512_ net26 VGND VGND VPWR VPWR complete_votes\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5729_ _2714_ tree_instances\[19\].u_tree.frame_id_out\[2\] tree_instances\[19\].u_tree.prediction_valid
+ VGND VGND VPWR VPWR _2774_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_17_264 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_79_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6475__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6404__RESET_B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_11_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_102_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_629 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_23_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_46 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3362__A _0732_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4060_ _1535_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_64_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_19_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4962_ _2217_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_47_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6701_ clknet_leaf_63_clk _0097_ net35 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_44 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_74_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3913_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1393_ sky130_fd_sc_hd__inv_2
X_4893_ _0953_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[7\] VGND
+ VGND VPWR VPWR _2173_ sky130_fd_sc_hd__or2_1
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6632_ clknet_leaf_64_clk _0391_ net35 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_197 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3844_ _1328_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3775_ _1264_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__clkbuf_1
X_6563_ clknet_leaf_18_clk _0081_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_54_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_595 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6986__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6494_ clknet_leaf_101_clk _0277_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[3\]
+ sky130_fd_sc_hd__dfxtp_1
X_5514_ net7 _0000_ _2574_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_42_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5445_ tree_instances\[1\].u_tree.tree_state\[1\] _0865_ _1820_ VGND VGND VPWR VPWR
+ _2533_ sky130_fd_sc_hd__or3_1
XANTENNA__6915__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_626 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_66_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5376_ _2465_ VGND VGND VPWR VPWR _2478_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4368__A _1112_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_74_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_484 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4327_ _1793_ VGND VGND VPWR VPWR _1794_ sky130_fd_sc_hd__clkbuf_1
X_4258_ _1696_ VGND VGND VPWR VPWR _1727_ sky130_fd_sc_hd__clkbuf_1
X_3209_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[7\] _0758_ VGND VGND
+ VPWR VPWR _0759_ sky130_fd_sc_hd__nor2_1
X_4189_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _1661_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_429 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_80_616 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5708__A2 _2600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6656__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3182__A _0733_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_EDGE_ROW_16_Right_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_16_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_44_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3560_ tree_instances\[14\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_25_Right_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6397__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3491_ _1001_ _1008_ _1017_ tree_instances\[7\].u_tree.tree_state\[1\] VGND VGND
+ VPWR VPWR _0082_ sky130_fd_sc_hd__a31o_1
X_5230_ tree_instances\[17\].u_tree.frame_id_out\[2\] tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0909_ VGND VGND VPWR VPWR _2386_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_110_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6326__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5161_ _2334_ VGND VGND VPWR VPWR _2335_ sky130_fd_sc_hd__clkbuf_1
X_5092_ tree_instances\[16\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _2290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4112_ _1165_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__clkbuf_1
X_4043_ _1511_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_3_Left_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_34_Right_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_108_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_108_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5994_ _2956_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__clkbuf_1
X_4945_ _1721_ _2133_ VGND VGND VPWR VPWR _2209_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_602 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5747__A _2586_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_454 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_19_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4876_ _2156_ VGND VGND VPWR VPWR _2157_ sky130_fd_sc_hd__clkbuf_1
X_6615_ clknet_leaf_50_clk _0378_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_valid\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_EDGE_ROW_43_Right_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3827_ tree_instances\[10\].u_tree.prediction_valid _1136_ VGND VGND VPWR VPWR _1315_
+ sky130_fd_sc_hd__and2b_1
X_6546_ clknet_leaf_44_clk _0320_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3758_ _0732_ tree_instances\[19\].u_tree.pipeline_valid\[0\] VGND VGND VPWR VPWR
+ _1251_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_76_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6477_ clknet_leaf_10_clk _0265_ net25 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3689_ _1190_ _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__nand2_1
X_5428_ _2522_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5359_ _2455_ VGND VGND VPWR VPWR _2461_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_292 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_52_Right_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_524 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_281 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_41_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_67_Left_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_61_Right_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_638 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6837__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_589 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__3177__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_21_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_98_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_76_Left_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_EDGE_ROW_70_Right_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5617__A1 _2603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_49_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_57_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_29_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_85_Left_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5567__A _2579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4730_ _2059_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6578__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4661_ _2015_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3612_ tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[2\] VGND VGND VPWR
+ VPWR _1126_ sky130_fd_sc_hd__clkbuf_1
X_6400_ clknet_leaf_49_clk _0202_ net35 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4592_ _1970_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6865__SET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6507__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6331_ clknet_leaf_90_clk _0139_ net27 VGND VGND VPWR VPWR tree_instances\[8\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3543_ _1061_ _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3474_ tree_instances\[7\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__clkbuf_1
X_6262_ _3130_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__clkbuf_1
X_6193_ _1891_ _3035_ VGND VGND VPWR VPWR _3092_ sky130_fd_sc_hd__and2_1
X_5213_ _2377_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5856__A1 _1829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5144_ _2320_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_71_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5608__A1 _2600_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5608__B2 _2588_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5075_ _2281_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__clkbuf_1
X_4026_ _1502_ VGND VGND VPWR VPWR _1503_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6033__A1 _0799_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5977_ _1329_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[3\] tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[4\]
+ _1319_ VGND VGND VPWR VPWR _2944_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_82_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4595__A1 _1835_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4928_ _1718_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[7\] _2192_
+ VGND VGND VPWR VPWR _2200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6930__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_7_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_573 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4859_ _0825_ VGND VGND VPWR VPWR _2140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_351 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_6529_ clknet_leaf_37_clk _0079_ net30 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_253 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_100_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_82_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_4
XTAP_TAPCELL_ROW_54_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6671__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6600__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_343 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_0_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3190_ tree_instances\[18\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _0743_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6263__A1 tree_instances\[0\].u_tree.frame_id_in\[4\] VGND VGND VPWR VPWR
+ sky130_fd_sc_hd__diode_2
XFILLER_0_72_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5900_ _2896_ VGND VGND VPWR VPWR _2899_ sky130_fd_sc_hd__buf_2
XTAP_TAPCELL_ROW_105_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_EDGE_ROW_93_Left_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_365 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_72_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_73_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6880_ clknet_leaf_12_clk _0599_ net29 VGND VGND VPWR VPWR tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5831_ tree_instances\[1\].u_tree.tree_state\[1\] tree_instances\[1\].u_tree.current_node_data\[12\]
+ tree_instances\[1\].u_tree.node_data\[12\] _2549_ VGND VGND VPWR VPWR _2854_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_410 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6759__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5762_ tree_instances\[6\].u_tree.frame_id_out\[4\] VGND VGND VPWR VPWR _2807_ sky130_fd_sc_hd__inv_2
XFILLER_0_29_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_593 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4713_ _2047_ VGND VGND VPWR VPWR _2048_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5526__A0 _2583_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5693_ _2580_ _2730_ _2731_ _2737_ VGND VGND VPWR VPWR _2738_ sky130_fd_sc_hd__o211a_1
X_4644_ _1578_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[0\] tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[7\]
+ _1596_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__a22o_1
XANTENNA__6341__RESET_B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5744__B _2579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4575_ _1788_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[3\] _1956_
+ VGND VGND VPWR VPWR _1961_ sky130_fd_sc_hd__mux2_1
X_6314_ clknet_leaf_30_clk _0123_ net28 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3526_ _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__clkbuf_1
X_6245_ tree_instances\[5\].u_tree.u_tree_weight_rom.cached_addr\[5\] _2477_ _3116_
+ VGND VGND VPWR VPWR _3122_ sky130_fd_sc_hd__mux2_1
X_3457_ _0980_ _0986_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__nand2_1
XANTENNA__5760__A _2659_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3388_ tree_instances\[16\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _0925_ sky130_fd_sc_hd__buf_1
X_6176_ tree_instances\[5\].u_tree.tree_state\[0\] tree_instances\[5\].u_tree.tree_state\[1\]
+ tree_instances\[5\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _3083_ sky130_fd_sc_hd__nor3_1
X_5127_ tree_instances\[16\].u_tree.read_enable VGND VGND VPWR VPWR _2310_ sky130_fd_sc_hd__inv_2
X_5058_ _2272_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__clkbuf_1
XPHY_EDGE_ROW_2_Right_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4009_ _1486_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_84_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_64_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA__6006__A1 _1829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_109_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_35_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_101_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_59_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_630 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_3_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_55_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6852__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_161 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_100_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_449 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5564__B _2613_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4360_ _1112_ tree_instances\[9\].u_tree.pipeline_valid\[0\] tree_instances\[9\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_1_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3311_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__clkbuf_1
X_4291_ _1758_ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__clkbuf_1
X_3242_ _0790_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__clkbuf_1
X_6030_ _2977_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__clkbuf_1
X_3173_ tree_instances\[4\].u_tree.tree_state\[2\] VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_46_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6932_ clknet_leaf_2_clk _0644_ VGND VGND VPWR VPWR tree_instances\[13\].u_tree.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_65_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6593__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6863_ clknet_leaf_85_clk _0583_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_TAPCELL_ROW_37_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5814_ _2845_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4362__C net1 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6794_ clknet_leaf_1_clk _0051_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.tree_state\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_29_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_390 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5745_ _2580_ tree_instances\[11\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2790_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5676_ tree_instances\[4\].u_tree.frame_id_out\[0\] VGND VGND VPWR VPWR _2721_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4627_ tree_instances\[9\].u_tree.tree_state\[0\] _1024_ VGND VGND VPWR VPWR _1988_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_25_490 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_102_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4558_ _1755_ _1945_ VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__and2_1
XTAP_TAPCELL_ROW_9_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4489_ _1791_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[1\] _1910_
+ _1036_ VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__o22a_1
X_3509_ _0846_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__clkbuf_1
X_6228_ _2361_ VGND VGND VPWR VPWR _3111_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_90_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_90_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5683__C1 _2727_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6159_ _2959_ VGND VGND VPWR VPWR _3068_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_37_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_644 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_79_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_67_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_29 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_90_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput5 net5 VGND VGND VPWR VPWR frame_id_out[3] sky130_fd_sc_hd__buf_8
XANTENNA_clkbuf_leaf_94_clk_A clknet_3_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_28_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_102_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_62_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_58_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_34_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3860_ _1317_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__clkbuf_1
X_3791_ _1280_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_32_clk_A clknet_3_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5530_ _2586_ net5 _1020_ VGND VGND VPWR VPWR _2587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_14_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5461_ _1498_ _2533_ VGND VGND VPWR VPWR _2542_ sky130_fd_sc_hd__and2_1
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4412_ tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1846_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_47_clk_A clknet_3_6__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5392_ tree_instances\[8\].u_tree.pipeline_valid\[0\] tree_instances\[8\].u_tree.tree_state\[0\]
+ VGND VGND VPWR VPWR _2494_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_EDGE_ROW_99_Right_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4343_ _1805_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__buf_2
X_4274_ _1741_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_6_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3225_ _0757_ _0761_ _0770_ _0774_ tree_instances\[20\].u_tree.tree_state\[1\] VGND
+ VGND VPWR VPWR _0070_ sky130_fd_sc_hd__a41o_1
X_6013_ _2966_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__clkbuf_1
X_3156_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_70 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6774__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_68_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_19_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_4
XANTENNA__6703__RESET_B net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6915_ clknet_leaf_31_clk _0628_ net29 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.frame_id_out\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_49_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6846_ clknet_leaf_66_clk _0566_ tree_instances\[0\].u_tree.rst_n VGND VGND VPWR
+ VPWR tree_instances\[2\].u_tree.pipeline_frame_id\[0\]\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_407 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_91_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6777_ clknet_leaf_6_clk _0511_ net26 VGND VGND VPWR VPWR complete_votes\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3989_ _1467_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__clkbuf_1
X_5728_ _2709_ tree_instances\[19\].u_tree.frame_id_out\[3\] _2772_ _2589_ VGND VGND
+ VPWR VPWR _2773_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_79_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5659_ _2573_ _0000_ VGND VGND VPWR VPWR _2705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_102_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_471 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6444__RESET_B net24 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_11_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_27 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_59_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_19_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4961_ tree_instances\[12\].u_tree.current_node_data\[12\] tree_instances\[12\].u_tree.node_data\[12\]
+ _1026_ VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_47_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6700_ clknet_leaf_55_clk _0449_ net37 VGND VGND VPWR VPWR tree_instances\[19\].u_tree.ready_for_next
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_80_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3912_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1392_ sky130_fd_sc_hd__clkbuf_1
X_4892_ _0953_ tree_instances\[13\].u_tree.u_tree_weight_rom.cached_addr\[7\] VGND
+ VGND VPWR VPWR _2172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6631_ clknet_leaf_64_clk _0390_ net35 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.pipeline_frame_id\[0\]\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3843_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[3\] VGND VGND VPWR
+ VPWR _1328_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_96 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3774_ _1263_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__clkbuf_1
X_6562_ clknet_leaf_44_clk _0092_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_319 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_54_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6493_ clknet_leaf_101_clk _0276_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[2\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5513_ _2571_ _2572_ _0000_ _2573_ VGND VGND VPWR VPWR _2574_ sky130_fd_sc_hd__o211a_1
X_5444_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_data\[12\] _2529_ _2532_
+ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_8_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5375_ _2476_ VGND VGND VPWR VPWR _2477_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_74_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_496 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4326_ _1049_ VGND VGND VPWR VPWR _1793_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6955__RESET_B tree_instances\[0\].u_tree.rst_n VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4257_ _1725_ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6752__SET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3208_ tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _0758_ sky130_fd_sc_hd__buf_1
X_4188_ tree_instances\[13\].u_tree.pipeline_current_node\[0\]\[5\] VGND VGND VPWR
+ VPWR _1660_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6829_ clknet_leaf_39_clk _0550_ net30 VGND VGND VPWR VPWR tree_instances\[1\].u_tree.frame_id_out\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3728__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_628 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_393 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_60_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6696__RESET_B net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_3 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6625__RESET_B net38 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_39 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_49 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_68_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_16_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_TAPCELL_ROW_44_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_max_cap27_A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_50_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6014__A _0032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_544 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3490_ _1012_ _1016_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_110_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5160_ _2333_ VGND VGND VPWR VPWR _2334_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6366__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5091_ _1137_ _2289_ _2275_ tree_instances\[15\].u_tree.ready_for_next VGND VGND
+ VPWR VPWR _0354_ sky130_fd_sc_hd__a22o_1
X_4111_ _1575_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__clkbuf_1
X_4042_ _1517_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_108_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5993_ tree_instances\[20\].u_tree.u_tree_weight_rom.cached_addr\[3\] _1432_ _2899_
+ VGND VGND VPWR VPWR _2956_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_474 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4944_ _2208_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4875_ _0818_ VGND VGND VPWR VPWR _2156_ sky130_fd_sc_hd__clkbuf_1
X_6614_ clknet_leaf_38_clk _0094_ net30 VGND VGND VPWR VPWR tree_instances\[16\].u_tree.prediction_valid
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3826_ _1314_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_168 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_104_218 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XPHY_EDGE_ROW_104_Left_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6545_ clknet_leaf_44_clk _0319_ net34 VGND VGND VPWR VPWR tree_instances\[14\].u_tree.pipeline_frame_id\[0\]\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_15_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3757_ _1245_ _1246_ _1250_ tree_instances\[5\].u_tree.tree_state\[2\] VGND VGND
+ VPWR VPWR _0035_ sky130_fd_sc_hd__o31a_1
XANTENNA__5571__A1 _2619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_76_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_588 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6476_ clknet_leaf_100_clk _0264_ net26 VGND VGND VPWR VPWR tree_instances\[12\].u_tree.read_enable
+ sky130_fd_sc_hd__dfrtp_2
X_3688_ _1191_ _1192_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__nor2_1
X_5427_ _1494_ tree_instances\[1\].u_tree.u_tree_weight_rom.cached_addr\[2\] _2519_
+ VGND VGND VPWR VPWR _2522_ sky130_fd_sc_hd__mux2_1
X_5358_ tree_instances\[5\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _2460_ sky130_fd_sc_hd__inv_2
X_4309_ tree_instances\[8\].u_tree.pipeline_current_node\[0\]\[1\] VGND VGND VPWR
+ VPWR _1776_ sky130_fd_sc_hd__inv_2
X_5289_ tree_instances\[18\].u_tree.frame_id_out\[2\] tree_instances\[18\].u_tree.pipeline_frame_id\[0\]\[2\]
+ _0753_ VGND VGND VPWR VPWR _2417_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_536 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_87_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_41_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_308 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_18_382 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5562__A1 _2585_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_98_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_21_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6806__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_49_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_45_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_29_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_57_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4660_ _1638_ _2012_ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_477 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_9_15 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3611_ tree_instances\[0\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1125_ sky130_fd_sc_hd__clkbuf_1
X_6330_ clknet_leaf_21_clk _0138_ net24 VGND VGND VPWR VPWR tree_instances\[7\].u_tree.pipeline_current_node\[0\]\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4591_ tree_instances\[9\].u_tree.pipeline_frame_id\[0\]\[1\] _1830_ _0044_ VGND
+ VGND VPWR VPWR _1970_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_650 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_12_503 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3542_ _1062_ tree_instances\[15\].u_tree.pipeline_current_node\[0\]\[4\] VGND VGND
+ VPWR VPWR _1063_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_246 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_86_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6261_ tree_instances\[6\].u_tree.pipeline_frame_id\[0\]\[3\] _1834_ _0038_ VGND
+ VGND VPWR VPWR _3130_ sky130_fd_sc_hd__mux2_1
X_3473_ tree_instances\[8\].u_tree.tree_state\[0\] _0999_ _1000_ VGND VGND VPWR VPWR
+ _0083_ sky130_fd_sc_hd__a21o_1
XANTENNA__6547__RESET_B net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6192_ _3091_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__clkbuf_1
X_5212_ _2376_ _2366_ VGND VGND VPWR VPWR _2377_ sky130_fd_sc_hd__and2_1
X_5143_ tree_instances\[16\].u_tree.prediction_out tree_instances\[16\].u_tree.pipeline_prediction\[0\]\[0\]
+ tree_instances\[16\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _2320_ sky130_fd_sc_hd__mux2_1
XTAP_TAPCELL_ROW_71_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5522__S _1020_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5074_ _1534_ _2255_ VGND VGND VPWR VPWR _2281_ sky130_fd_sc_hd__and2_1
X_4025_ tree_instances\[19\].u_tree.pipeline_current_node\[0\]\[0\] VGND VGND VPWR
+ VPWR _1502_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5758__A _2622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_219 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5976_ _1189_ _2939_ _2940_ _2942_ VGND VGND VPWR VPWR _2943_ sky130_fd_sc_hd__a211o_1
XTAP_TAPCELL_ROW_82_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4927_ _2199_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_425 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_7_541 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4858_ _0829_ _0830_ _1810_ tree_instances\[12\].u_tree.ready_for_next VGND VGND
+ VPWR VPWR _0271_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3809_ _1288_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_585 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_34_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4789_ _1702_ tree_instances\[12\].u_tree.u_tree_weight_rom.cached_addr\[0\] _2091_
+ _0839_ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6528_ clknet_leaf_59_clk _0062_ net38 VGND VGND VPWR VPWR tree_instances\[17\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_6459_ clknet_leaf_24_clk _0034_ net24 VGND VGND VPWR VPWR tree_instances\[4\].u_tree.tree_state\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_265 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__5668__A _2603_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_54_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_26_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_455 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_108_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__6640__RESET_B net35 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_355 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_333 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_88_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_105_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5830_ _1934_ tree_instances\[8\].u_tree.node_data\[12\] _2853_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_data\[12\]
+ _1967_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_422 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5761_ _2603_ tree_instances\[6\].u_tree.frame_id_out\[1\] tree_instances\[6\].u_tree.frame_id_out\[4\]
+ _2708_ _2805_ VGND VGND VPWR VPWR _2806_ sky130_fd_sc_hd__o221a_1
X_4712_ _2046_ VGND VGND VPWR VPWR _2047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_617 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XANTENNA__6799__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5692_ _2734_ _2735_ _2736_ VGND VGND VPWR VPWR _2737_ sky130_fd_sc_hd__nor3_1
XFILLER_0_56_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4643_ _1579_ tree_instances\[10\].u_tree.u_tree_weight_rom.cached_addr\[0\] _2000_
+ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_533 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_4_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6728__RESET_B net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4574_ _1960_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_94 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6313_ clknet_leaf_30_clk _0122_ net28 VGND VGND VPWR VPWR tree_instances\[6\].u_tree.pipeline_current_node\[0\]\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_3525_ _1046_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6381__RESET_B net39 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6244_ _3121_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__6310__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3456_ _0983_ _0985_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__nor2_1
X_3387_ _0923_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__clkbuf_1
X_6175_ tree_instances\[5\].u_tree.tree_state\[1\] tree_instances\[5\].u_tree.current_node_data\[107\]
+ tree_instances\[5\].u_tree.node_data\[107\] _0933_ VGND VGND VPWR VPWR _3082_ sky130_fd_sc_hd__a22o_1
X_5126_ _2309_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__clkbuf_1
X_5057_ tree_instances\[15\].u_tree.pipeline_frame_id\[0\]\[2\] _2125_ _0016_ VGND
+ VGND VPWR VPWR _2272_ sky130_fd_sc_hd__mux2_1
X_4008_ _1476_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__clkbuf_1
XTAP_TAPCELL_ROW_84_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_84_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_51_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_23_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5959_ _1418_ _2552_ VGND VGND VPWR VPWR _2930_ sky130_fd_sc_hd__and2_1
XFILLER_0_75_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_47_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6469__RESET_B net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_105_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_95_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_30_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3471__A _0731_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_59_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_98_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_TAPCELL_ROW_3_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_641 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_53_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_173 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XTAP_TAPCELL_ROW_100_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6821__RESET_B net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_130 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_349 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3310_ tree_instances\[3\].u_tree.pipeline_current_node\[0\]\[5\] _0852_ VGND VGND
+ VPWR VPWR _0853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4290_ _1745_ VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_174 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3241_ tree_instances\[17\].u_tree.pipeline_current_node\[0\]\[6\] VGND VGND VPWR
+ VPWR _0790_ sky130_fd_sc_hd__inv_2
XFILLER_0_67_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3172_ _0722_ _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_6_clk_A clknet_3_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6931_ clknet_leaf_100_clk _0643_ VGND VGND VPWR VPWR tree_instances\[12\].u_tree.node_data\[12\]
+ sky130_fd_sc_hd__dfxtp_1
XFILLER_0_49_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6862_ clknet_leaf_76_clk _0582_ net39 VGND VGND VPWR VPWR tree_instances\[20\].u_tree.pipeline_current_node\[0\]\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5813_ tree_instances\[0\].u_tree.pipeline_frame_id\[0\]\[3\] _2249_ _0004_ VGND
+ VGND VPWR VPWR _2845_ sky130_fd_sc_hd__mux2_1
X_6793_ clknet_leaf_48_clk _0046_ net34 VGND VGND VPWR VPWR tree_instances\[0\].u_tree.tree_state\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__6909__RESET_B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5744_ tree_instances\[11\].u_tree.frame_id_out\[1\] _2579_ VGND VGND VPWR VPWR _2789_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_17_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6562__RESET_B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5675_ _2580_ tree_instances\[4\].u_tree.frame_id_out\[1\] VGND VGND VPWR VPWR _2720_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4626_ _1987_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4557_ _1951_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4488_ tree_instances\[8\].u_tree.u_tree_weight_rom.cached_addr\[6\] VGND VGND VPWR
+ VPWR _1910_ sky130_fd_sc_hd__inv_2
X_3508_ tree_instances\[12\].u_tree.pipeline_current_node\[0\]\[7\] VGND VGND VPWR
+ VPWR _1031_ sky130_fd_sc_hd__clkbuf_1
X_6227_ _2311_ VGND VGND VPWR VPWR _3110_ sky130_fd_sc_hd__clkbuf_1
X_3439_ tree_instances\[7\].u_tree.tree_state\[3\] VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__buf_2
XANTENNA__4387__A _1829_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_TAPCELL_ROW_90_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6158_ _1227_ _3067_ _0026_ tree_instances\[1\].u_tree.pipeline_valid\[0\] VGND VGND
+ VPWR VPWR _0645_ sky130_fd_sc_hd__o2bb2a_1
X_5109_ _1456_ _2296_ VGND VGND VPWR VPWR _2301_ sky130_fd_sc_hd__and2_1
XFILLER_0_57_90 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_6089_ tree_instances\[3\].u_tree.u_tree_weight_rom.cached_addr\[7\] _1346_ _3020_
+ VGND VGND VPWR VPWR _3024_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_TAPCELL_ROW_0_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_94_166 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_94_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput6 net6 VGND VGND VPWR VPWR frame_id_out[4] sky130_fd_sc_hd__buf_8
XFILLER_0_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_101_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_TAPCELL_ROW_102_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_85_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_TAPCELL_ROW_62_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_TAPCELL_ROW_34_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5729__A1 _2714_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_561 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_3790_ _1279_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_TAPCELL_ROW_14_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5460_ _2541_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_266 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4411_ _1845_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_225 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_41_247 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
XFILLER_0_10_601 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_5391_ _2491_ _2451_ _2488_ VGND VGND VPWR VPWR _2493_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_461 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4342_ tree_instances\[17\].u_tree.pipeline_valid\[0\] tree_instances\[17\].u_tree.tree_state\[0\]
+ net1 VGND VGND VPWR VPWR _1805_ sky130_fd_sc_hd__and3b_1
XFILLER_0_10_645 VPWR VGND VPWR VGND sky130_ef_sc_hd__decap_12
X_4273_ _1739_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__clkbuf_1
X_3224_ _0773_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__clkbuf_1
X_6012_ tree_instances\[3\].u_tree.pipeline_frame_id\[0\]\[4\] tree_instances\[0\].u_tree.frame_id_in\[4\]
+ _0032_ VGND VGND VPWR VPWR _2966_ sky130_fd_sc_hd__mux2_1
.ends

