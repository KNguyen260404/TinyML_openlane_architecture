module tree_rom_2 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000140681000000000000010023;
    rom[1] = 120'h001300000000000000000000001;
    rom[2] = 120'h0021407F3800000000000030883;
    rom[3] = 120'h00314077C800000000000040553;
    rom[4] = 120'h004041D8EC33500000000050343;
    rom[5] = 120'h005A40AEF800000000000060193;
    rom[6] = 120'h006A3FF000000000000000700E3;
    rom[7] = 120'h0071406890000000000000800B3;
    rom[8] = 120'h0081406830000000000000900A3;
    rom[9] = 120'h009300000000000000000000001;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B14068B0000000000000C00D3;
    rom[12] = 120'h00C300000000000000000000000;
    rom[13] = 120'h00D300000000000000000000001;
    rom[14] = 120'h00EA402900000000000000F0143;
    rom[15] = 120'h00FA40040000000000000100113;
    rom[16] = 120'h010300000000000000000000000;
    rom[17] = 120'h011A40240000000000000120133;
    rom[18] = 120'h012300000000000000000000001;
    rom[19] = 120'h013300000000000000000000000;
    rom[20] = 120'h0141406E3000000000000150183;
    rom[21] = 120'h015A40504000000000000160173;
    rom[22] = 120'h016300000000000000000000000;
    rom[23] = 120'h017300000000000000000000001;
    rom[24] = 120'h018300000000000000000000001;
    rom[25] = 120'h019A43D1C0F3A000000001A0293;
    rom[26] = 120'h01A1406F30000000000001B0223;
    rom[27] = 120'h01B1406930000000000001C01F3;
    rom[28] = 120'h01CA43CA7C732000000001D01E3;
    rom[29] = 120'h01D300000000000000000000000;
    rom[30] = 120'h01E300000000000000000000001;
    rom[31] = 120'h01F1406E1000000000000200213;
    rom[32] = 120'h020300000000000000000000001;
    rom[33] = 120'h021300000000000000000000000;
    rom[34] = 120'h022140734800000000000230263;
    rom[35] = 120'h023A43D19E79D00000000240253;
    rom[36] = 120'h024300000000000000000000001;
    rom[37] = 120'h025300000000000000000000000;
    rom[38] = 120'h026A4211FCE6000000000270283;
    rom[39] = 120'h027300000000000000000000001;
    rom[40] = 120'h028300000000000000000000001;
    rom[41] = 120'h0291406F30000000000002A02F3;
    rom[42] = 120'h02AA43DF7718D000000002B02E3;
    rom[43] = 120'h02BA43DEC150A000000002C02D3;
    rom[44] = 120'h02C300000000000000000000001;
    rom[45] = 120'h02D300000000000000000000000;
    rom[46] = 120'h02E300000000000000000000001;
    rom[47] = 120'h02FA43D5BBBD700000000300313;
    rom[48] = 120'h030300000000000000000000001;
    rom[49] = 120'h03114072A800000000000320333;
    rom[50] = 120'h032300000000000000000000001;
    rom[51] = 120'h033300000000000000000000001;
    rom[52] = 120'h034041D8EC33B00000000350543;
    rom[53] = 120'h035041D8EC33700000000360453;
    rom[54] = 120'h036A40AFDC000000000003703E3;
    rom[55] = 120'h03714068B0000000000003803B3;
    rom[56] = 120'h038A404C00000000000003903A3;
    rom[57] = 120'h039300000000000000000000000;
    rom[58] = 120'h03A300000000000000000000001;
    rom[59] = 120'h03BA402700000000000003C03D3;
    rom[60] = 120'h03C300000000000000000000001;
    rom[61] = 120'h03D300000000000000000000001;
    rom[62] = 120'h03EA43CA1A5CE000000003F0423;
    rom[63] = 120'h03F1406F3000000000000400413;
    rom[64] = 120'h040300000000000000000000000;
    rom[65] = 120'h041300000000000000000000001;
    rom[66] = 120'h042A43D1C6B7600000000430443;
    rom[67] = 120'h043300000000000000000000001;
    rom[68] = 120'h044300000000000000000000001;
    rom[69] = 120'h045A40A6B6000000000004604D3;
    rom[70] = 120'h0461407318000000000004704A3;
    rom[71] = 120'h047041D8EC33900000000480493;
    rom[72] = 120'h048300000000000000000000001;
    rom[73] = 120'h049300000000000000000000001;
    rom[74] = 120'h04A041D8EC339000000004B04C3;
    rom[75] = 120'h04B300000000000000000000001;
    rom[76] = 120'h04C300000000000000000000000;
    rom[77] = 120'h04DA43D206BA1000000004E0513;
    rom[78] = 120'h04E1407348000000000004F0503;
    rom[79] = 120'h04F300000000000000000000000;
    rom[80] = 120'h050300000000000000000000001;
    rom[81] = 120'h051041D8EC33900000000520533;
    rom[82] = 120'h052300000000000000000000001;
    rom[83] = 120'h053300000000000000000000000;
    rom[84] = 120'h054300000000000000000000000;
    rom[85] = 120'h055041D8EC33900000000560873;
    rom[86] = 120'h056041D8EC33700000000570703;
    rom[87] = 120'h057A43EA3A50A00000000580673;
    rom[88] = 120'h058041D8EC33500000000590603;
    rom[89] = 120'h0591407E58000000000005A05D3;
    rom[90] = 120'h05AA43D40CF61000000005B05C3;
    rom[91] = 120'h05B300000000000000000000000;
    rom[92] = 120'h05C300000000000000000000000;
    rom[93] = 120'h05D1407F08000000000005E05F3;
    rom[94] = 120'h05E300000000000000000000001;
    rom[95] = 120'h05F300000000000000000000000;
    rom[96] = 120'h0601407E5800000000000610643;
    rom[97] = 120'h0611407A1800000000000620633;
    rom[98] = 120'h062300000000000000000000000;
    rom[99] = 120'h063300000000000000000000000;
    rom[100] = 120'h064A43240018100000000650663;
    rom[101] = 120'h065300000000000000000000001;
    rom[102] = 120'h066300000000000000000000000;
    rom[103] = 120'h067A43EB0072B000000006806F3;
    rom[104] = 120'h068041D8EC335000000006906C3;
    rom[105] = 120'h06914079A8000000000006A06B3;
    rom[106] = 120'h06A300000000000000000000001;
    rom[107] = 120'h06B300000000000000000000001;
    rom[108] = 120'h06C14079B8000000000006D06E3;
    rom[109] = 120'h06D300000000000000000000001;
    rom[110] = 120'h06E300000000000000000000001;
    rom[111] = 120'h06F300000000000000000000001;
    rom[112] = 120'h0701407E60000000000007107A3;
    rom[113] = 120'h071A43EA163C600000000720793;
    rom[114] = 120'h072A43D44D36400000000730763;
    rom[115] = 120'h073A41EEBF0DA00000000740753;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h075300000000000000000000000;
    rom[118] = 120'h076A43DFDE11200000000770783;
    rom[119] = 120'h077300000000000000000000001;
    rom[120] = 120'h078300000000000000000000000;
    rom[121] = 120'h079300000000000000000000001;
    rom[122] = 120'h07AA432500180000000007B0823;
    rom[123] = 120'h07B1407F28000000000007C07F3;
    rom[124] = 120'h07C1407E98000000000007D07E3;
    rom[125] = 120'h07D300000000000000000000001;
    rom[126] = 120'h07E300000000000000000000001;
    rom[127] = 120'h07FA415119BDE00000000800813;
    rom[128] = 120'h080300000000000000000000000;
    rom[129] = 120'h081300000000000000000000001;
    rom[130] = 120'h082A43E6F906A00000000830863;
    rom[131] = 120'h0831407F1800000000000840853;
    rom[132] = 120'h084300000000000000000000000;
    rom[133] = 120'h085300000000000000000000001;
    rom[134] = 120'h086300000000000000000000001;
    rom[135] = 120'h087300000000000000000000000;
    rom[136] = 120'h088041D8EC33900000000890D63;
    rom[137] = 120'h089041D8EC337000000008A0B93;
    rom[138] = 120'h08AA3FE000000000000008B09C3;
    rom[139] = 120'h08B041D8EC335000000008C0953;
    rom[140] = 120'h08C14088D8000000000008D08E3;
    rom[141] = 120'h08D300000000000000000000001;
    rom[142] = 120'h08E1409002000000000008F0923;
    rom[143] = 120'h08F1408C5800000000000900913;
    rom[144] = 120'h090300000000000000000000000;
    rom[145] = 120'h091300000000000000000000000;
    rom[146] = 120'h09214092C000000000000930943;
    rom[147] = 120'h093300000000000000000000001;
    rom[148] = 120'h094300000000000000000000000;
    rom[149] = 120'h0951408930000000000001200973;
    rom[150] = 120'h0120300000000000000000000001;
    rom[151] = 120'h09714091AA00000000000980993;
    rom[152] = 120'h098300000000000000000000000;
    rom[153] = 120'h09914093B4000000000009A09B3;
    rom[154] = 120'h09A300000000000000000000001;
    rom[155] = 120'h09B300000000000000000000000;
    rom[156] = 120'h09C1408FDC000000000009D0AC3;
    rom[157] = 120'h09D1408F64000000000009E0A53;
    rom[158] = 120'h09EA43B2F2DFE000000009F0A23;
    rom[159] = 120'h09F041D8EC33500000000A00A13;
    rom[160] = 120'h0A0300000000000000000000001;
    rom[161] = 120'h0A1300000000000000000000001;
    rom[162] = 120'h0A21408F4400000000000A30A43;
    rom[163] = 120'h0A3300000000000000000000001;
    rom[164] = 120'h0A4300000000000000000000001;
    rom[165] = 120'h0A51408F6C00000000000A60A93;
    rom[166] = 120'h0A6A43DF0C73100000000A70A83;
    rom[167] = 120'h0A7300000000000000000000001;
    rom[168] = 120'h0A8300000000000000000000000;
    rom[169] = 120'h0A91408FC400000000000AA0AB3;
    rom[170] = 120'h0AA300000000000000000000001;
    rom[171] = 120'h0AB300000000000000000000000;
    rom[172] = 120'h0AC14094AA00000000000AD0B43;
    rom[173] = 120'h0AD041D8EC33500000000AE0B13;
    rom[174] = 120'h0AE140930200000000000AF0B03;
    rom[175] = 120'h0AF300000000000000000000001;
    rom[176] = 120'h0B0300000000000000000000001;
    rom[177] = 120'h0B1140930200000000000B20B33;
    rom[178] = 120'h0B2300000000000000000000001;
    rom[179] = 120'h0B3300000000000000000000001;
    rom[180] = 120'h0B4A42D0011EF00000000B50B83;
    rom[181] = 120'h0B51409DC200000000000B60B73;
    rom[182] = 120'h0B6300000000000000000000001;
    rom[183] = 120'h0B7300000000000000000000001;
    rom[184] = 120'h0B8300000000000000000000001;
    rom[185] = 120'h0B9140861400000000000BA0C73;
    rom[186] = 120'h0BAA43917FC4700000000BB0C03;
    rom[187] = 120'h0BB1407F5800000000000BC0BF3;
    rom[188] = 120'h0BCA43601000400FDFB40BD0BE3;
    rom[189] = 120'h0BD300000000000000000000001;
    rom[190] = 120'h0BE300000000000000000000000;
    rom[191] = 120'h0BF300000000000000000000001;
    rom[192] = 120'h0C01407F5800000000000C10C63;
    rom[193] = 120'h0C11407F4800000000000C20C33;
    rom[194] = 120'h0C2300000000000000000000001;
    rom[195] = 120'h0C3A43B90900100000000C40C53;
    rom[196] = 120'h0C4300000000000000000000001;
    rom[197] = 120'h0C5300000000000000000000000;
    rom[198] = 120'h0C6300000000000000000000001;
    rom[199] = 120'h0C7A3FE00000000000000C80C93;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C91408E8C00000000000CA0CF3;
    rom[202] = 120'h0CAA439F90EA600000000CB0CE3;
    rom[203] = 120'h0CB1408E0400000000000CC0CD3;
    rom[204] = 120'h0CC300000000000000000000000;
    rom[205] = 120'h0CD300000000000000000000000;
    rom[206] = 120'h0CE300000000000000000000001;
    rom[207] = 120'h0CFA426C1D38700000000D00D33;
    rom[208] = 120'h0D0A40840400000000000D10D23;
    rom[209] = 120'h0D1300000000000000000000001;
    rom[210] = 120'h0D2300000000000000000000001;
    rom[211] = 120'h0D31408F6400000000000D40D53;
    rom[212] = 120'h0D4300000000000000000000001;
    rom[213] = 120'h0D5300000000000000000000001;
    rom[214] = 120'h0D6041D8EC33B00000000D70E83;
    rom[215] = 120'h0D7A421EC808700000000D80E13;
    rom[216] = 120'h0D81408CCC00000000000D90DE3;
    rom[217] = 120'h0D91408A4800000000000DA0DB3;
    rom[218] = 120'h0DA300000000000000000000000;
    rom[219] = 120'h0DBA4201C1B515C000000DC0DD3;
    rom[220] = 120'h0DC300000000000000000000000;
    rom[221] = 120'h0DD300000000000000000000001;
    rom[222] = 120'h0DEA41E00000270000000DF0E03;
    rom[223] = 120'h0DF300000000000000000000000;
    rom[224] = 120'h0E0300000000000000000000001;
    rom[225] = 120'h0E114082E000000000000E20E73;
    rom[226] = 120'h0E2A43A13000080000000E30E43;
    rom[227] = 120'h0E3300000000000000000000000;
    rom[228] = 120'h0E4A43AB1B00000000000E50E63;
    rom[229] = 120'h0E5300000000000000000000001;
    rom[230] = 120'h0E6300000000000000000000000;
    rom[231] = 120'h0E7300000000000000000000000;
    rom[232] = 120'h0E81408EE800000000000E90EA3;
    rom[233] = 120'h0E9300000000000000000000000;
    rom[234] = 120'h0EA041D8EC33D00000000EB0F03;
    rom[235] = 120'h0EBA43BBF184C00000000EC0ED3;
    rom[236] = 120'h0EC300000000000000000000000;
    rom[237] = 120'h0EDA43C02A4F780000000EE0EF3;
    rom[238] = 120'h0EE300000000000000000000001;
    rom[239] = 120'h0EF300000000000000000000000;
    rom[240] = 120'h0F0041D8EC33F00000000F10F63;
    rom[241] = 120'h0F1A425D680B800000000F20F53;
    rom[242] = 120'h0F2A42140000040000000F30F43;
    rom[243] = 120'h0F3300000000000000000000000;
    rom[244] = 120'h0F4300000000000000000000001;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 

