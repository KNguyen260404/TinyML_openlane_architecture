module tree_rom_16 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000041D8EC339000000000112E3;
    rom[1] = 120'h001A43C2154BD00000000020CB3;
    rom[2] = 120'h002A4360009A700000000030663;
    rom[3] = 120'h003A432318AC300000000040373;
    rom[4] = 120'h0041406E10000000000000501A3;
    rom[5] = 120'h005A40CFD4000000000000600D3;
    rom[6] = 120'h006140681000000000000070083;
    rom[7] = 120'h007300000000000000000000001;
    rom[8] = 120'h00814068D0000000000000900C3;
    rom[9] = 120'h009041D8EC335000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000000;
    rom[12] = 120'h00C300000000000000000000001;
    rom[13] = 120'h00D041D8EC337000000000E0153;
    rom[14] = 120'h00EA40D04D200000000000F0123;
    rom[15] = 120'h00F1406A6000000000000100113;
    rom[16] = 120'h010300000000000000000000000;
    rom[17] = 120'h011300000000000000000000001;
    rom[18] = 120'h012140681000000000000130143;
    rom[19] = 120'h013300000000000000000000001;
    rom[20] = 120'h014300000000000000000000001;
    rom[21] = 120'h015A42F40D62800000000160173;
    rom[22] = 120'h016300000000000000000000001;
    rom[23] = 120'h017140692000000000000180193;
    rom[24] = 120'h018300000000000000000000000;
    rom[25] = 120'h019300000000000000000000001;
    rom[26] = 120'h01A041D8EC337000000001B02A3;
    rom[27] = 120'h01B041D8EC335000000001C0233;
    rom[28] = 120'h01CA3FE000000000000001D0203;
    rom[29] = 120'h01D1409002000000000001E01F3;
    rom[30] = 120'h01E300000000000000000000000;
    rom[31] = 120'h01F300000000000000000000000;
    rom[32] = 120'h0201407E9800000000000210223;
    rom[33] = 120'h021300000000000000000000000;
    rom[34] = 120'h022300000000000000000000001;
    rom[35] = 120'h0231408A5400000000000240273;
    rom[36] = 120'h024A3FF00000000000000250263;
    rom[37] = 120'h025300000000000000000000000;
    rom[38] = 120'h026300000000000000000000000;
    rom[39] = 120'h027A3FE00000000000000280293;
    rom[40] = 120'h028300000000000000000000000;
    rom[41] = 120'h029300000000000000000000001;
    rom[42] = 120'h02A1408A5C000000000002B0303;
    rom[43] = 120'h02BA3FF000000000000002C02D3;
    rom[44] = 120'h02C300000000000000000000000;
    rom[45] = 120'h02D1407E98000000000002E02F3;
    rom[46] = 120'h02E300000000000000000000000;
    rom[47] = 120'h02F300000000000000000000000;
    rom[48] = 120'h0301408FCC00000000000310343;
    rom[49] = 120'h0311408F4400000000000320333;
    rom[50] = 120'h032300000000000000000000001;
    rom[51] = 120'h033300000000000000000000001;
    rom[52] = 120'h034A400C0000000000000350363;
    rom[53] = 120'h035300000000000000000000000;
    rom[54] = 120'h036300000000000000000000001;
    rom[55] = 120'h037041D8EC335000000003804B3;
    rom[56] = 120'h038A4324356C6000000003903C3;
    rom[57] = 120'h0391407550000000000003A03B3;
    rom[58] = 120'h03A300000000000000000000000;
    rom[59] = 120'h03B300000000000000000000001;
    rom[60] = 120'h03CA43528175D000000003D0443;
    rom[61] = 120'h03DA4351DDDCB000000003E0413;
    rom[62] = 120'h03EA434384C88000000003F0403;
    rom[63] = 120'h03F300000000000000000000001;
    rom[64] = 120'h040300000000000000000000001;
    rom[65] = 120'h041A4351E5A1F00000000420433;
    rom[66] = 120'h042300000000000000000000000;
    rom[67] = 120'h043300000000000000000000001;
    rom[68] = 120'h044140692000000000000450483;
    rom[69] = 120'h045140681000000000000460473;
    rom[70] = 120'h046300000000000000000000001;
    rom[71] = 120'h047300000000000000000000000;
    rom[72] = 120'h048A435B7D71E000000004904A3;
    rom[73] = 120'h049300000000000000000000001;
    rom[74] = 120'h04A300000000000000000000001;
    rom[75] = 120'h04BA4329F9344000000004C0573;
    rom[76] = 120'h04C1407028000000000004D0503;
    rom[77] = 120'h04D14067B0000000000004E04F3;
    rom[78] = 120'h04E300000000000000000000001;
    rom[79] = 120'h04F300000000000000000000000;
    rom[80] = 120'h050A43240018100000000510543;
    rom[81] = 120'h051041D8EC33700000000520533;
    rom[82] = 120'h052300000000000000000000001;
    rom[83] = 120'h053300000000000000000000001;
    rom[84] = 120'h054041D8EC33700000000550563;
    rom[85] = 120'h055300000000000000000000001;
    rom[86] = 120'h056300000000000000000000001;
    rom[87] = 120'h05714068D0000000000005805F3;
    rom[88] = 120'h058A433E8F021000000005905C3;
    rom[89] = 120'h059A433D9FB59000000005A05B3;
    rom[90] = 120'h05A300000000000000000000000;
    rom[91] = 120'h05B300000000000000000000001;
    rom[92] = 120'h05C1406810000000000005D05E3;
    rom[93] = 120'h05D300000000000000000000001;
    rom[94] = 120'h05E300000000000000000000000;
    rom[95] = 120'h05FA4354B151400000000600633;
    rom[96] = 120'h060A43468B7B200000000610623;
    rom[97] = 120'h061300000000000000000000001;
    rom[98] = 120'h062300000000000000000000001;
    rom[99] = 120'h0631407E7000000000000640653;
    rom[100] = 120'h064300000000000000000000001;
    rom[101] = 120'h065300000000000000000000001;
    rom[102] = 120'h066041D8EC33700000000670A43;
    rom[103] = 120'h0671407E9800000000000680873;
    rom[104] = 120'h068A437002BB100000000690783;
    rom[105] = 120'h069041D8EC335000000006A0713;
    rom[106] = 120'h06AA436089840000000006B06E3;
    rom[107] = 120'h06B14069D0000000000006C06D3;
    rom[108] = 120'h06C300000000000000000000000;
    rom[109] = 120'h06D300000000000000000000001;
    rom[110] = 120'h06EA436EC661C000000006F0703;
    rom[111] = 120'h06F300000000000000000000001;
    rom[112] = 120'h070300000000000000000000000;
    rom[113] = 120'h071A4360815FC00000000720753;
    rom[114] = 120'h072A436014CFE00000000730743;
    rom[115] = 120'h073300000000000000000000000;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h075A43666308100000000760773;
    rom[118] = 120'h076300000000000000000000001;
    rom[119] = 120'h077300000000000000000000000;
    rom[120] = 120'h078A43B0E066D00000000790803;
    rom[121] = 120'h079041D8EC335000000007A07D3;
    rom[122] = 120'h07AA43A001DE7000000007B07C3;
    rom[123] = 120'h07B300000000000000000000000;
    rom[124] = 120'h07C300000000000000000000000;
    rom[125] = 120'h07DA43A13D1CF000000007E07F3;
    rom[126] = 120'h07E300000000000000000000000;
    rom[127] = 120'h07F300000000000000000000000;
    rom[128] = 120'h08014068B000000000000810843;
    rom[129] = 120'h081041D8EC33500000000820833;
    rom[130] = 120'h082300000000000000000000000;
    rom[131] = 120'h083300000000000000000000000;
    rom[132] = 120'h084041D8EC33500000000850863;
    rom[133] = 120'h085300000000000000000000001;
    rom[134] = 120'h086300000000000000000000001;
    rom[135] = 120'h087041D8EC33500000000880953;
    rom[136] = 120'h0881407F70000000000008908E3;
    rom[137] = 120'h089A43AF91C82000000008A08D3;
    rom[138] = 120'h08A1407F48000000000008B08C3;
    rom[139] = 120'h08B300000000000000000000001;
    rom[140] = 120'h08C300000000000000000000000;
    rom[141] = 120'h08D300000000000000000000001;
    rom[142] = 120'h08E1408F8C000000000008F0923;
    rom[143] = 120'h08FA439EE351D00000000900913;
    rom[144] = 120'h090300000000000000000000000;
    rom[145] = 120'h091300000000000000000000001;
    rom[146] = 120'h09214094AC00000000000930943;
    rom[147] = 120'h093300000000000000000000001;
    rom[148] = 120'h094300000000000000000000001;
    rom[149] = 120'h095A43A000E41000000009609D3;
    rom[150] = 120'h096A4374B0000000000009709A3;
    rom[151] = 120'h0971407F7000000000000980993;
    rom[152] = 120'h098300000000000000000000000;
    rom[153] = 120'h099300000000000000000000001;
    rom[154] = 120'h09A1408F6C000000000009B09C3;
    rom[155] = 120'h09B300000000000000000000000;
    rom[156] = 120'h09C300000000000000000000001;
    rom[157] = 120'h09DA43AB9695A000000009E0A13;
    rom[158] = 120'h09E1408F20000000000009F0A03;
    rom[159] = 120'h09F300000000000000000000001;
    rom[160] = 120'h0A0300000000000000000000001;
    rom[161] = 120'h0A1A43AE1E00200000000A20A33;
    rom[162] = 120'h0A2300000000000000000000000;
    rom[163] = 120'h0A3300000000000000000000001;
    rom[164] = 120'h0A4A43A1A484C00000000A50B63;
    rom[165] = 120'h0A514093F600000000000A60B53;
    rom[166] = 120'h0A6A436FF2FB100000000A70AE3;
    rom[167] = 120'h0A7140706800000000000A80AB3;
    rom[168] = 120'h0A8A43600600200000000A90AA3;
    rom[169] = 120'h0A9300000000000000000000000;
    rom[170] = 120'h0AA300000000000000000000000;
    rom[171] = 120'h0AB1408F4000000000000AC0AD3;
    rom[172] = 120'h0AC300000000000000000000001;
    rom[173] = 120'h0AD300000000000000000000000;
    rom[174] = 120'h0AEA43A0C48AB00000000AF0B23;
    rom[175] = 120'h0AF140631000000000000B00B13;
    rom[176] = 120'h0B0300000000000000000000001;
    rom[177] = 120'h0B1300000000000000000000000;
    rom[178] = 120'h0B21408CF400000000000B30B43;
    rom[179] = 120'h0B3300000000000000000000001;
    rom[180] = 120'h0B4300000000000000000000000;
    rom[181] = 120'h0B5300000000000000000000001;
    rom[182] = 120'h0B61407E9800000000000B70BE3;
    rom[183] = 120'h0B7140673000000000000B80B93;
    rom[184] = 120'h0B8300000000000000000000001;
    rom[185] = 120'h0B9A43AC7F17400000000BA0BB3;
    rom[186] = 120'h0BA300000000000000000000001;
    rom[187] = 120'h0BB140695000000000000BC0BD3;
    rom[188] = 120'h0BC300000000000000000000000;
    rom[189] = 120'h0BD300000000000000000000000;
    rom[190] = 120'h0BE140930000000000000BF0C63;
    rom[191] = 120'h0BF1408F3400000000000C00C33;
    rom[192] = 120'h0C0A43C1D376D00000000C10C23;
    rom[193] = 120'h0C1300000000000000000000001;
    rom[194] = 120'h0C2300000000000000000000000;
    rom[195] = 120'h0C3A43B33A1C400000000C40C53;
    rom[196] = 120'h0C4300000000000000000000000;
    rom[197] = 120'h0C5300000000000000000000001;
    rom[198] = 120'h0C614094B800000000000C70CA3;
    rom[199] = 120'h0C714094A200000000000C80C93;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C9300000000000000000000000;
    rom[202] = 120'h0CA300000000000000000000001;
    rom[203] = 120'h0CB041D8EC33700000000CC1033;
    rom[204] = 120'h0CCA43C7FFB4800000000CD0CE3;
    rom[205] = 120'h0CD300000000000000000000001;
    rom[206] = 120'h0CE041D8EC33500000000CF0EA3;
    rom[207] = 120'h0CFA43D3FFF6000000000D00DD3;
    rom[208] = 120'h0D01407E9800000000000D10D83;
    rom[209] = 120'h0D1A43D17BFC600000000D20D53;
    rom[210] = 120'h0D2A43D00C49D00000000D30D43;
    rom[211] = 120'h0D3300000000000000000000000;
    rom[212] = 120'h0D4300000000000000000000001;
    rom[213] = 120'h0D5A43D1C0F3A00000000D60D73;
    rom[214] = 120'h0D6300000000000000000000000;
    rom[215] = 120'h0D7300000000000000000000000;
    rom[216] = 120'h0D8140932200000000000D90DA3;
    rom[217] = 120'h0D9300000000000000000000001;
    rom[218] = 120'h0DA140932600000000000DB0DC3;
    rom[219] = 120'h0DB300000000000000000000000;
    rom[220] = 120'h0DC300000000000000000000001;
    rom[221] = 120'h0DD1407F1800000000000DE0E53;
    rom[222] = 120'h0DE140798800000000000DF0E23;
    rom[223] = 120'h0DFA43DED7D4B00000000E00E13;
    rom[224] = 120'h0E0300000000000000000000001;
    rom[225] = 120'h0E1300000000000000000000001;
    rom[226] = 120'h0E2A43EA3BB6300000000E30E43;
    rom[227] = 120'h0E3300000000000000000000000;
    rom[228] = 120'h0E4300000000000000000000001;
    rom[229] = 120'h0E51408F6C00000000000E60E93;
    rom[230] = 120'h0E61408F6400000000000E70E83;
    rom[231] = 120'h0E7300000000000000000000001;
    rom[232] = 120'h0E8300000000000000000000000;
    rom[233] = 120'h0E9300000000000000000000001;
    rom[234] = 120'h0EA1407F1800000000000EB0FA3;
    rom[235] = 120'h0EB140798800000000000EC0F33;
    rom[236] = 120'h0ECA43CA14FBE00000000ED0F03;
    rom[237] = 120'h0EDA43C88860F00000000EE0EF3;
    rom[238] = 120'h0EE300000000000000000000000;
    rom[239] = 120'h0EF300000000000000000000000;
    rom[240] = 120'h0F0140729800000000000F10F23;
    rom[241] = 120'h0F1300000000000000000000001;
    rom[242] = 120'h0F2300000000000000000000001;
    rom[243] = 120'h0F314079D800000000000F40F73;
    rom[244] = 120'h0F4A43EB4F93600000000F50F63;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
