module tree_rom_12 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000A43C2154C500000000010E83;
    rom[1] = 120'h001041D8EC33900000000020B53;
    rom[2] = 120'h002041D8EC33500000000030443;
    rom[3] = 120'h003140689000000000000040133;
    rom[4] = 120'h004140681000000000000050063;
    rom[5] = 120'h005300000000000000000000001;
    rom[6] = 120'h006140683000000000000070123;
    rom[7] = 120'h007A4203FB67E000000000800B3;
    rom[8] = 120'h008A403700000000000000900A3;
    rom[9] = 120'h009300000000000000000000001;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00BA42DFA87E5000000000C00F3;
    rom[12] = 120'h00CA4255E46D0300000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00FA43A8E3C2400000000100113;
    rom[16] = 120'h010300000000000000000000000;
    rom[17] = 120'h011300000000000000000000000;
    rom[18] = 120'h012300000000000000000000001;
    rom[19] = 120'h013A3FE00000000000000140253;
    rom[20] = 120'h0141409002000000000001501E3;
    rom[21] = 120'h015140726000000000000160193;
    rom[22] = 120'h016140692000000000000170183;
    rom[23] = 120'h017300000000000000000000000;
    rom[24] = 120'h018300000000000000000000001;
    rom[25] = 120'h0191408014000000000001A01B3;
    rom[26] = 120'h01A300000000000000000000000;
    rom[27] = 120'h01B14088D8000000000001C01D3;
    rom[28] = 120'h01C300000000000000000000001;
    rom[29] = 120'h01D300000000000000000000000;
    rom[30] = 120'h01E14092C0000000000001F0203;
    rom[31] = 120'h01F300000000000000000000001;
    rom[32] = 120'h0201409D0600000000000210243;
    rom[33] = 120'h021140950C00000000000220233;
    rom[34] = 120'h022300000000000000000000000;
    rom[35] = 120'h023300000000000000000000001;
    rom[36] = 120'h024300000000000000000000000;
    rom[37] = 120'h025A417007B4E00000000260353;
    rom[38] = 120'h026A4138BC1A0000000002702E3;
    rom[39] = 120'h0271407E18000000000002802B3;
    rom[40] = 120'h0281407E08000000000002902A3;
    rom[41] = 120'h029300000000000000000000001;
    rom[42] = 120'h02A300000000000000000000000;
    rom[43] = 120'h02BA408038000000000002C02D3;
    rom[44] = 120'h02C300000000000000000000001;
    rom[45] = 120'h02D300000000000000000000001;
    rom[46] = 120'h02EA416D9F70B000000002F0323;
    rom[47] = 120'h02FA41629EA5300000000300313;
    rom[48] = 120'h030300000000000000000000001;
    rom[49] = 120'h031300000000000000000000001;
    rom[50] = 120'h032A416DA08A300000000330343;
    rom[51] = 120'h033300000000000000000000000;
    rom[52] = 120'h034300000000000000000000001;
    rom[53] = 120'h035A436FEB0F4000000003603D3;
    rom[54] = 120'h0361407E18000000000003703A3;
    rom[55] = 120'h037A41EF934BC00000000380393;
    rom[56] = 120'h038300000000000000000000000;
    rom[57] = 120'h039300000000000000000000000;
    rom[58] = 120'h03AA4196FC49B000000003B03C3;
    rom[59] = 120'h03B300000000000000000000000;
    rom[60] = 120'h03C300000000000000000000001;
    rom[61] = 120'h03D1407F58000000000003E0413;
    rom[62] = 120'h03EA43B230D49000000003F0403;
    rom[63] = 120'h03F300000000000000000000000;
    rom[64] = 120'h040300000000000000000000000;
    rom[65] = 120'h041A439DA30AF00000000420433;
    rom[66] = 120'h042300000000000000000000000;
    rom[67] = 120'h043300000000000000000000001;
    rom[68] = 120'h044041D8EC33700000000450803;
    rom[69] = 120'h0451408A5400000000000460653;
    rom[70] = 120'h046A436000A0A00000000470563;
    rom[71] = 120'h047A432023627000000004804F3;
    rom[72] = 120'h048A417071201000000004904C3;
    rom[73] = 120'h049A400400000000000004A04B3;
    rom[74] = 120'h04A300000000000000000000000;
    rom[75] = 120'h04B300000000000000000000001;
    rom[76] = 120'h04C1406810000000000004D04E3;
    rom[77] = 120'h04D300000000000000000000001;
    rom[78] = 120'h04E300000000000000000000000;
    rom[79] = 120'h04FA43240018100000000500533;
    rom[80] = 120'h0501406C4000000000000510523;
    rom[81] = 120'h051300000000000000000000001;
    rom[82] = 120'h052300000000000000000000001;
    rom[83] = 120'h053A435F49A9A00000000540553;
    rom[84] = 120'h054300000000000000000000001;
    rom[85] = 120'h055300000000000000000000001;
    rom[86] = 120'h056A43A1182AA000000005705E3;
    rom[87] = 120'h057A437002BB1000000005805B3;
    rom[88] = 120'h058A4360815FC000000005905A3;
    rom[89] = 120'h059300000000000000000000000;
    rom[90] = 120'h05A300000000000000000000001;
    rom[91] = 120'h05BA439925C4A000000005C05D3;
    rom[92] = 120'h05C300000000000000000000000;
    rom[93] = 120'h05D300000000000000000000000;
    rom[94] = 120'h05EA43AE09AC5000000005F0623;
    rom[95] = 120'h05F1407E9800000000000600613;
    rom[96] = 120'h060300000000000000000000001;
    rom[97] = 120'h061300000000000000000000001;
    rom[98] = 120'h0621407F7000000000000630643;
    rom[99] = 120'h063300000000000000000000000;
    rom[100] = 120'h064300000000000000000000001;
    rom[101] = 120'h0651408FDC00000000000660753;
    rom[102] = 120'h066A4374B0000000000006706E3;
    rom[103] = 120'h0671408F84000000000006806B3;
    rom[104] = 120'h0681408E84000000000006906A3;
    rom[105] = 120'h069300000000000000000000001;
    rom[106] = 120'h06A300000000000000000000001;
    rom[107] = 120'h06BA430AA0048800000006C06D3;
    rom[108] = 120'h06C300000000000000000000000;
    rom[109] = 120'h06D300000000000000000000000;
    rom[110] = 120'h06EA43B3381C4000000006F0723;
    rom[111] = 120'h06FA439F288E000000000700713;
    rom[112] = 120'h070300000000000000000000000;
    rom[113] = 120'h071300000000000000000000000;
    rom[114] = 120'h072A43B79E7FA00000000730743;
    rom[115] = 120'h073300000000000000000000001;
    rom[116] = 120'h074300000000000000000000001;
    rom[117] = 120'h075A3FE000000000000007607B3;
    rom[118] = 120'h07614093B400000000000770783;
    rom[119] = 120'h077300000000000000000000001;
    rom[120] = 120'h07814099A6000000000007907A3;
    rom[121] = 120'h079300000000000000000000000;
    rom[122] = 120'h07A300000000000000000000000;
    rom[123] = 120'h07BA43C20A073000000007C07F3;
    rom[124] = 120'h07C14093C6000000000007D07E3;
    rom[125] = 120'h07D300000000000000000000001;
    rom[126] = 120'h07E300000000000000000000001;
    rom[127] = 120'h07F300000000000000000000000;
    rom[128] = 120'h080A43A0C47D9000000008109C3;
    rom[129] = 120'h0811408E8C000000000008208F3;
    rom[130] = 120'h082A435F9DD77000000008308A3;
    rom[131] = 120'h083A43224626500000000840873;
    rom[132] = 120'h0841406E1000000000000850863;
    rom[133] = 120'h085300000000000000000000001;
    rom[134] = 120'h086300000000000000000000000;
    rom[135] = 120'h087A4329C74E000000000880893;
    rom[136] = 120'h088300000000000000000000001;
    rom[137] = 120'h089300000000000000000000000;
    rom[138] = 120'h08A1406800000000000008B08C3;
    rom[139] = 120'h08B300000000000000000000001;
    rom[140] = 120'h08CA43666F018000000008D08E3;
    rom[141] = 120'h08D300000000000000000000000;
    rom[142] = 120'h08E300000000000000000000000;
    rom[143] = 120'h08FA426C1D38700000000900953;
    rom[144] = 120'h0901408FCC00000000000910923;
    rom[145] = 120'h091300000000000000000000001;
    rom[146] = 120'h092A40840400000000000930943;
    rom[147] = 120'h093300000000000000000000000;
    rom[148] = 120'h094300000000000000000000001;
    rom[149] = 120'h0951408FD800000000000960993;
    rom[150] = 120'h096A4337AFBA400000000970983;
    rom[151] = 120'h097300000000000000000000000;
    rom[152] = 120'h098300000000000000000000000;
    rom[153] = 120'h09914093C6000000000009A09B3;
    rom[154] = 120'h09A300000000000000000000001;
    rom[155] = 120'h09B300000000000000000000001;
    rom[156] = 120'h09CA43AE930A5000000009D0A63;
    rom[157] = 120'h09D1408F30000000000009E0A33;
    rom[158] = 120'h09E1407ED8000000000009F0A23;
    rom[159] = 120'h09F1407D7800000000000A00A13;
    rom[160] = 120'h0A0300000000000000000000001;
    rom[161] = 120'h0A1300000000000000000000000;
    rom[162] = 120'h0A2300000000000000000000001;
    rom[163] = 120'h0A31408FA400000000000A40A53;
    rom[164] = 120'h0A4300000000000000000000000;
    rom[165] = 120'h0A5300000000000000000000001;
    rom[166] = 120'h0A6A43B33C50E00000000A70AE3;
    rom[167] = 120'h0A7A43AF2F8F800000000A80AB3;
    rom[168] = 120'h0A81408F6800000000000A90AA3;
    rom[169] = 120'h0A9300000000000000000000000;
    rom[170] = 120'h0AA300000000000000000000001;
    rom[171] = 120'h0AB140930C00000000000AC0AD3;
    rom[172] = 120'h0AC300000000000000000000000;
    rom[173] = 120'h0AD300000000000000000000001;
    rom[174] = 120'h0AE14068B000000000000AF0B23;
    rom[175] = 120'h0AFA43C20656600000000B00B13;
    rom[176] = 120'h0B0300000000000000000000000;
    rom[177] = 120'h0B1300000000000000000000001;
    rom[178] = 120'h0B214094A200000000000B30B43;
    rom[179] = 120'h0B3300000000000000000000001;
    rom[180] = 120'h0B4300000000000000000000001;
    rom[181] = 120'h0B5041D8EC33B00000000B60D73;
    rom[182] = 120'h0B6A42D00000200000000B70CE3;
    rom[183] = 120'h0B71406BA000000000000B80BF3;
    rom[184] = 120'h0B8A419C0082100000000B90BE3;
    rom[185] = 120'h0B9A40C00800000000000BA0BB3;
    rom[186] = 120'h0BA300000000000000000000001;
    rom[187] = 120'h0BBA418C0104200000000BC0BD3;
    rom[188] = 120'h0BC300000000000000000000000;
    rom[189] = 120'h0BD300000000000000000000001;
    rom[190] = 120'h0BE300000000000000000000000;
    rom[191] = 120'h0BFA41EFF150000000000C00C53;
    rom[192] = 120'h0C0A41300104800000000C10C23;
    rom[193] = 120'h0C1300000000000000000000000;
    rom[194] = 120'h0C2A41300A0F800000000C30C43;
    rom[195] = 120'h0C3300000000000000000000001;
    rom[196] = 120'h0C4300000000000000000000000;
    rom[197] = 120'h0C5140890C00000000000C60C93;
    rom[198] = 120'h0C614073E800000000000C70C83;
    rom[199] = 120'h0C7300000000000000000000001;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C9140917400000000000CA0CD3;
    rom[202] = 120'h0CAA42654630838000000CB0CC3;
    rom[203] = 120'h0CB300000000000000000000001;
    rom[204] = 120'h0CC300000000000000000000000;
    rom[205] = 120'h0CD300000000000000000000000;
    rom[206] = 120'h0CEA43AA0919500000000CF0D03;
    rom[207] = 120'h0CF300000000000000000000000;
    rom[208] = 120'h0D01407EF000000000000D10D23;
    rom[209] = 120'h0D1300000000000000000000000;
    rom[210] = 120'h0D2140877800000000000D30D63;
    rom[211] = 120'h0D3A43AB1B00000000000D40D53;
    rom[212] = 120'h0D4300000000000000000000001;
    rom[213] = 120'h0D5300000000000000000000000;
    rom[214] = 120'h0D6300000000000000000000000;
    rom[215] = 120'h0D7041D8EC33D00000000D80DF3;
    rom[216] = 120'h0D81408EE800000000000D90DA3;
    rom[217] = 120'h0D9300000000000000000000000;
    rom[218] = 120'h0DA1408F6800000000000DB0DE3;
    rom[219] = 120'h0DBA43BBF184C00000000DC0DD3;
    rom[220] = 120'h0DC300000000000000000000000;
    rom[221] = 120'h0DD300000000000000000000001;
    rom[222] = 120'h0DE300000000000000000000000;
    rom[223] = 120'h0DF041D8EC33F00000000E00E73;
    rom[224] = 120'h0E01408EE800000000000E10E23;
    rom[225] = 120'h0E1300000000000000000000000;
    rom[226] = 120'h0E2A425D680B800000000E30E63;
    rom[227] = 120'h0E3A42140000040000000E40E53;
    rom[228] = 120'h0E4300000000000000000000000;
    rom[229] = 120'h0E5300000000000000000000001;
    rom[230] = 120'h0E6300000000000000000000000;
    rom[231] = 120'h0E7300000000000000000000000;
    rom[232] = 120'h0E8140681000000000000E90EA3;
    rom[233] = 120'h0E9300000000000000000000001;
    rom[234] = 120'h0EA1407F5800000000000EB1283;
    rom[235] = 120'h0EBA43D3FFF6000000000EC1033;
    rom[236] = 120'h0EC1407E9800000000000ED0FA3;
    rom[237] = 120'h0EDA43C7FFB4800000000EE0EF3;
    rom[238] = 120'h0EE300000000000000000000001;
    rom[239] = 120'h0EF140798800000000000F00F53;
    rom[240] = 120'h0F0041D8EC33900000000F10F43;
    rom[241] = 120'h0F114068B000000000000F20F33;
    rom[242] = 120'h0F2300000000000000000000000;
    rom[243] = 120'h0F3300000000000000000000001;
    rom[244] = 120'h0F4300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
