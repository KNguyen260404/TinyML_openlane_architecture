module tree_rom_19 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000A43C2154C500000000010FE3;
    rom[1] = 120'h001A43600000C000000000207B3;
    rom[2] = 120'h0021406E1000000000000030283;
    rom[3] = 120'h003041D8EC33B00000000040273;
    rom[4] = 120'h004140689000000000000050143;
    rom[5] = 120'h005A42F03F535800000000600F3;
    rom[6] = 120'h006140681000000000000070083;
    rom[7] = 120'h007300000000000000000000001;
    rom[8] = 120'h008A4203FB67E000000000900C3;
    rom[9] = 120'h0091406830000000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00C1406830000000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00F140681000000000000100113;
    rom[16] = 120'h010300000000000000000000001;
    rom[17] = 120'h011140683000000000000120133;
    rom[18] = 120'h012300000000000000000000000;
    rom[19] = 120'h013300000000000000000000001;
    rom[20] = 120'h014A40CED280000000000150183;
    rom[21] = 120'h01514068C000000000000160173;
    rom[22] = 120'h016300000000000000000000000;
    rom[23] = 120'h017300000000000000000000001;
    rom[24] = 120'h018041D8EC33500000000190203;
    rom[25] = 120'h019A41AB463A6000000001A01D3;
    rom[26] = 120'h01AA419A143C2000000001B01C3;
    rom[27] = 120'h01B300000000000000000000001;
    rom[28] = 120'h01C300000000000000000000000;
    rom[29] = 120'h01D14068B0000000000001E01F3;
    rom[30] = 120'h01E300000000000000000000000;
    rom[31] = 120'h01F300000000000000000000001;
    rom[32] = 120'h020041D8EC33900000000210243;
    rom[33] = 120'h02114068B000000000000220233;
    rom[34] = 120'h022300000000000000000000000;
    rom[35] = 120'h023300000000000000000000001;
    rom[36] = 120'h02414068E000000000000250263;
    rom[37] = 120'h025300000000000000000000000;
    rom[38] = 120'h026300000000000000000000001;
    rom[39] = 120'h027300000000000000000000000;
    rom[40] = 120'h0281408A5400000000000290563;
    rom[41] = 120'h029041D8EC339000000002A0493;
    rom[42] = 120'h02A041D8EC337000000002B03A3;
    rom[43] = 120'h02B1407E18000000000002C0333;
    rom[44] = 120'h02C041D8EC335000000002D0303;
    rom[45] = 120'h02D1406F30000000000002E02F3;
    rom[46] = 120'h02E300000000000000000000000;
    rom[47] = 120'h02F300000000000000000000000;
    rom[48] = 120'h030A431C6016900000000310323;
    rom[49] = 120'h031300000000000000000000000;
    rom[50] = 120'h032300000000000000000000001;
    rom[51] = 120'h033A3FE00000000000000340373;
    rom[52] = 120'h034140893000000000000350363;
    rom[53] = 120'h035300000000000000000000000;
    rom[54] = 120'h036300000000000000000000000;
    rom[55] = 120'h037041D8EC33500000000380393;
    rom[56] = 120'h038300000000000000000000001;
    rom[57] = 120'h039300000000000000000000001;
    rom[58] = 120'h03A1407E18000000000003B0423;
    rom[59] = 120'h03B14077E8000000000003C03F3;
    rom[60] = 120'h03C1407388000000000003D03E3;
    rom[61] = 120'h03D300000000000000000000000;
    rom[62] = 120'h03E300000000000000000000001;
    rom[63] = 120'h03F1407CD800000000000400413;
    rom[64] = 120'h040300000000000000000000000;
    rom[65] = 120'h041300000000000000000000000;
    rom[66] = 120'h0421407F2800000000000430463;
    rom[67] = 120'h0431407E9800000000000440453;
    rom[68] = 120'h044300000000000000000000001;
    rom[69] = 120'h045300000000000000000000001;
    rom[70] = 120'h046A42A5CECDD00000000470483;
    rom[71] = 120'h047300000000000000000000000;
    rom[72] = 120'h048300000000000000000000001;
    rom[73] = 120'h04914075F8000000000004A0513;
    rom[74] = 120'h04A1406EA0000000000004B04C3;
    rom[75] = 120'h04B300000000000000000000000;
    rom[76] = 120'h04C041D8EC33B000000004D0503;
    rom[77] = 120'h04DA412012090000000004E04F3;
    rom[78] = 120'h04E300000000000000000000000;
    rom[79] = 120'h04F300000000000000000000001;
    rom[80] = 120'h050300000000000000000000000;
    rom[81] = 120'h0511408A4800000000000520533;
    rom[82] = 120'h052300000000000000000000000;
    rom[83] = 120'h053A4201C3DD180000000540553;
    rom[84] = 120'h054300000000000000000000000;
    rom[85] = 120'h055300000000000000000000001;
    rom[86] = 120'h0561409DC2000000000005706C3;
    rom[87] = 120'h057A3FE000000000000005805F3;
    rom[88] = 120'h058041D8EC337000000005905E3;
    rom[89] = 120'h0591409436000000000005A05D3;
    rom[90] = 120'h05A041D8EC335000000005B05C3;
    rom[91] = 120'h05B300000000000000000000000;
    rom[92] = 120'h05C300000000000000000000000;
    rom[93] = 120'h05D300000000000000000000001;
    rom[94] = 120'h05E300000000000000000000000;
    rom[95] = 120'h05F041D8EC33B00000000600673;
    rom[96] = 120'h060041D8EC33900000000610643;
    rom[97] = 120'h061041D8EC33700000000620633;
    rom[98] = 120'h062300000000000000000000001;
    rom[99] = 120'h063300000000000000000000001;
    rom[100] = 120'h064A425C480B800000000650663;
    rom[101] = 120'h065300000000000000000000001;
    rom[102] = 120'h066300000000000000000000000;
    rom[103] = 120'h067A425D680B8000000006806B3;
    rom[104] = 120'h068A4214000004E0000006906A3;
    rom[105] = 120'h069300000000000000000000000;
    rom[106] = 120'h06A300000000000000000000001;
    rom[107] = 120'h06B300000000000000000000000;
    rom[108] = 120'h06C041D8EC339000000006D07A3;
    rom[109] = 120'h06D1409DCE000000000006E0753;
    rom[110] = 120'h06E041D8EC335000000006F0723;
    rom[111] = 120'h06F1409DCA00000000000700713;
    rom[112] = 120'h070300000000000000000000000;
    rom[113] = 120'h071300000000000000000000000;
    rom[114] = 120'h072041D8EC33700000000730743;
    rom[115] = 120'h073300000000000000000000000;
    rom[116] = 120'h074300000000000000000000000;
    rom[117] = 120'h0751409DFE00000000000760793;
    rom[118] = 120'h076041D8EC33700000000770783;
    rom[119] = 120'h077300000000000000000000001;
    rom[120] = 120'h078300000000000000000000000;
    rom[121] = 120'h079300000000000000000000001;
    rom[122] = 120'h07A300000000000000000000000;
    rom[123] = 120'h07BA43A0B44F8000000007C0BF3;
    rom[124] = 120'h07CA4374B09A1000000007D0A43;
    rom[125] = 120'h07D1407F68000000000007E08D3;
    rom[126] = 120'h07EA436007208000000007F0843;
    rom[127] = 120'h07F14072D800000000000800813;
    rom[128] = 120'h080300000000000000000000000;
    rom[129] = 120'h081A436001A2700000000820833;
    rom[130] = 120'h082300000000000000000000000;
    rom[131] = 120'h083300000000000000000000001;
    rom[132] = 120'h084140680000000000000850863;
    rom[133] = 120'h085300000000000000000000001;
    rom[134] = 120'h0861406EE0000000000008708A3;
    rom[135] = 120'h087041D8EC33900000000880893;
    rom[136] = 120'h088300000000000000000000000;
    rom[137] = 120'h089300000000000000000000000;
    rom[138] = 120'h08AA43663B732000000008B08C3;
    rom[139] = 120'h08B300000000000000000000001;
    rom[140] = 120'h08C300000000000000000000000;
    rom[141] = 120'h08D1408FCC000000000008E09D3;
    rom[142] = 120'h08E041D8EC337000000008F0963;
    rom[143] = 120'h08FA4374A000000000000900933;
    rom[144] = 120'h090A436FE82AC00000000910923;
    rom[145] = 120'h091300000000000000000000001;
    rom[146] = 120'h092300000000000000000000000;
    rom[147] = 120'h093041D8EC33500000000940953;
    rom[148] = 120'h094300000000000000000000000;
    rom[149] = 120'h095300000000000000000000001;
    rom[150] = 120'h096A436989FF6000000009709A3;
    rom[151] = 120'h097041D8EC33900000000980993;
    rom[152] = 120'h098300000000000000000000001;
    rom[153] = 120'h099300000000000000000000000;
    rom[154] = 120'h09A041D8EC339000000009B09C3;
    rom[155] = 120'h09B300000000000000000000000;
    rom[156] = 120'h09C300000000000000000000000;
    rom[157] = 120'h09D041D8EC33B000000009E0A33;
    rom[158] = 120'h09E1409308000000000009F0A23;
    rom[159] = 120'h09F140930200000000000A00A13;
    rom[160] = 120'h0A0300000000000000000000001;
    rom[161] = 120'h0A1300000000000000000000000;
    rom[162] = 120'h0A2300000000000000000000001;
    rom[163] = 120'h0A3300000000000000000000000;
    rom[164] = 120'h0A414093C800000000000A50BE3;
    rom[165] = 120'h0A5A4399DB49B00000000A60B33;
    rom[166] = 120'h0A61407F6000000000000A70AE3;
    rom[167] = 120'h0A7041D8EC33700000000A80AB3;
    rom[168] = 120'h0A814067E000000000000A90AA3;
    rom[169] = 120'h0A9300000000000000000000001;
    rom[170] = 120'h0AA300000000000000000000000;
    rom[171] = 120'h0AB140639000000000000AC0AD3;
    rom[172] = 120'h0AC300000000000000000000001;
    rom[173] = 120'h0AD300000000000000000000000;
    rom[174] = 120'h0AE1408E7C00000000000AF0B03;
    rom[175] = 120'h0AF300000000000000000000001;
    rom[176] = 120'h0B0041D8EC33700000000B10B23;
    rom[177] = 120'h0B1300000000000000000000000;
    rom[178] = 120'h0B2300000000000000000000000;
    rom[179] = 120'h0B314078E800000000000B40B73;
    rom[180] = 120'h0B4041D8EC33900000000B50B63;
    rom[181] = 120'h0B5300000000000000000000001;
    rom[182] = 120'h0B6300000000000000000000000;
    rom[183] = 120'h0B7041D8EC33700000000B80BB3;
    rom[184] = 120'h0B8041D8EC33500000000B90BA3;
    rom[185] = 120'h0B9300000000000000000000000;
    rom[186] = 120'h0BA300000000000000000000000;
    rom[187] = 120'h0BBA439B1DD0800000000BC0BD3;
    rom[188] = 120'h0BC300000000000000000000000;
    rom[189] = 120'h0BD300000000000000000000000;
    rom[190] = 120'h0BE300000000000000000000001;
    rom[191] = 120'h0BF1407E9800000000000C00DD3;
    rom[192] = 120'h0C0140681000000000000C10C23;
    rom[193] = 120'h0C1300000000000000000000001;
    rom[194] = 120'h0C2041D8EC33700000000C30D23;
    rom[195] = 120'h0C314068B000000000000C40CB3;
    rom[196] = 120'h0C4041D8EC33500000000C50C83;
    rom[197] = 120'h0C5140689000000000000C60C73;
    rom[198] = 120'h0C6300000000000000000000000;
    rom[199] = 120'h0C7300000000000000000000000;
    rom[200] = 120'h0C8140689000000000000C90CA3;
    rom[201] = 120'h0C9300000000000000000000000;
    rom[202] = 120'h0CA300000000000000000000000;
    rom[203] = 120'h0CB041D8EC33500000000CC0CF3;
    rom[204] = 120'h0CC140798800000000000CD0CE3;
    rom[205] = 120'h0CD300000000000000000000001;
    rom[206] = 120'h0CE300000000000000000000000;
    rom[207] = 120'h0CFA43B009CF100000000D00D13;
    rom[208] = 120'h0D0300000000000000000000000;
    rom[209] = 120'h0D1300000000000000000000001;
    rom[210] = 120'h0D214068B000000000000D30D83;
    rom[211] = 120'h0D3A43BA750E200000000D40D73;
    rom[212] = 120'h0D4041D8EC33900000000D50D63;
    rom[213] = 120'h0D5300000000000000000000000;
    rom[214] = 120'h0D6300000000000000000000000;
    rom[215] = 120'h0D7300000000000000000000000;
    rom[216] = 120'h0D814078E800000000000D90DA3;
    rom[217] = 120'h0D9300000000000000000000001;
    rom[218] = 120'h0DAA43B37066D00000000DB0DC3;
    rom[219] = 120'h0DB300000000000000000000000;
    rom[220] = 120'h0DC300000000000000000000001;
    rom[221] = 120'h0DD041D8EC33900000000DE0F33;
    rom[222] = 120'h0DE1408F4000000000000DF0E83;
    rom[223] = 120'h0DF1407F5800000000000E00E73;
    rom[224] = 120'h0E0041D8EC33500000000E10E43;
    rom[225] = 120'h0E1A43AF91C8200000000E20E33;
    rom[226] = 120'h0E2300000000000000000000000;
    rom[227] = 120'h0E3300000000000000000000001;
    rom[228] = 120'h0E4A43C035FDD00000000E50E63;
    rom[229] = 120'h0E5300000000000000000000001;
    rom[230] = 120'h0E6300000000000000000000000;
    rom[231] = 120'h0E7300000000000000000000001;
    rom[232] = 120'h0E8041D8EC33500000000E90EE3;
    rom[233] = 120'h0E91408F4C00000000000EA0EB3;
    rom[234] = 120'h0EA300000000000000000000000;
    rom[235] = 120'h0EBA43C20FEBF00000000EC0ED3;
    rom[236] = 120'h0EC300000000000000000000001;
    rom[237] = 120'h0ED300000000000000000000000;
    rom[238] = 120'h0EE14094AA00000000000EF0F23;
    rom[239] = 120'h0EFA43B33B1C200000000F00F13;
    rom[240] = 120'h0F0300000000000000000000000;
    rom[241] = 120'h0F1300000000000000000000001;
    rom[242] = 120'h0F2300000000000000000000001;
    rom[243] = 120'h0F3A43AA1B17F00000000F40F73;
    rom[244] = 120'h0F4140877800000000000F50F63;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
