module Random_forest_top_ver2 (clk,
    feature_valid,
    prediction_out,
    prediction_valid,
    ready_for_next,
    rst_n,
    arbitration_id,
    data_field,
    frame_id_out,
    timestamp);
 input clk;
 input feature_valid;
 output prediction_out;
 output prediction_valid;
 output ready_for_next;
 input rst_n;
 input [63:0] arbitration_id;
 input [63:0] data_field;
 output [4:0] frame_id_out;
 input [63:0] timestamp;

 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire \attack_votes[0] ;
 wire \attack_votes[1] ;
 wire \attack_votes[2] ;
 wire \attack_votes[3] ;
 wire \attack_votes[4] ;
 wire \complete_votes[0] ;
 wire \complete_votes[1] ;
 wire \complete_votes[2] ;
 wire \complete_votes[3] ;
 wire \complete_votes[4] ;
 wire \current_voting_frame[0] ;
 wire \current_voting_frame[1] ;
 wire \current_voting_frame[2] ;
 wire \current_voting_frame[3] ;
 wire \current_voting_frame[4] ;
 wire \state[0] ;
 wire \state[1] ;
 wire \tree_instances[0].u_tree.frame_id_in[0] ;
 wire \tree_instances[0].u_tree.frame_id_in[1] ;
 wire \tree_instances[0].u_tree.frame_id_in[2] ;
 wire \tree_instances[0].u_tree.frame_id_in[3] ;
 wire \tree_instances[0].u_tree.frame_id_in[4] ;
 wire \tree_instances[0].u_tree.frame_id_out[0] ;
 wire \tree_instances[0].u_tree.frame_id_out[1] ;
 wire \tree_instances[0].u_tree.frame_id_out[2] ;
 wire \tree_instances[0].u_tree.frame_id_out[3] ;
 wire \tree_instances[0].u_tree.frame_id_out[4] ;
 wire \tree_instances[0].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[0].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[0].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[0].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[0].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[0].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[0].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[0].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[0].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[0].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[0].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[0].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[0].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[0].u_tree.pipeline_valid[0] ;
 wire \tree_instances[0].u_tree.prediction_valid ;
 wire \tree_instances[0].u_tree.ready_for_next ;
 wire \tree_instances[0].u_tree.rst_n ;
 wire \tree_instances[0].u_tree.tree_state[0] ;
 wire \tree_instances[0].u_tree.tree_state[1] ;
 wire \tree_instances[0].u_tree.tree_state[2] ;
 wire \tree_instances[0].u_tree.tree_state[3] ;
 wire \tree_instances[10].u_tree.current_node_data[12] ;
 wire \tree_instances[10].u_tree.frame_id_out[0] ;
 wire \tree_instances[10].u_tree.frame_id_out[1] ;
 wire \tree_instances[10].u_tree.frame_id_out[2] ;
 wire \tree_instances[10].u_tree.frame_id_out[3] ;
 wire \tree_instances[10].u_tree.frame_id_out[4] ;
 wire \tree_instances[10].u_tree.node_data[12] ;
 wire \tree_instances[10].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[10].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[10].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[10].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[10].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[10].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[10].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[10].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[10].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[10].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[10].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[10].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[10].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[10].u_tree.pipeline_prediction[0][0] ;
 wire \tree_instances[10].u_tree.pipeline_valid[0] ;
 wire \tree_instances[10].u_tree.prediction_out ;
 wire \tree_instances[10].u_tree.prediction_valid ;
 wire \tree_instances[10].u_tree.read_enable ;
 wire \tree_instances[10].u_tree.ready_for_next ;
 wire \tree_instances[10].u_tree.tree_state[0] ;
 wire \tree_instances[10].u_tree.tree_state[1] ;
 wire \tree_instances[10].u_tree.tree_state[2] ;
 wire \tree_instances[10].u_tree.tree_state[3] ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.cache_valid ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[0] ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[1] ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[2] ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[3] ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[4] ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[5] ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[6] ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[7] ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.cached_data[12] ;
 wire \tree_instances[10].u_tree.u_tree_weight_rom.gen_tree_10.u_tree_rom.node_data[12] ;
 wire \tree_instances[11].u_tree.frame_id_out[0] ;
 wire \tree_instances[11].u_tree.frame_id_out[1] ;
 wire \tree_instances[11].u_tree.frame_id_out[2] ;
 wire \tree_instances[11].u_tree.frame_id_out[3] ;
 wire \tree_instances[11].u_tree.frame_id_out[4] ;
 wire \tree_instances[11].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[11].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[11].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[11].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[11].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[11].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[11].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[11].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[11].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[11].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[11].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[11].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[11].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[11].u_tree.pipeline_valid[0] ;
 wire \tree_instances[11].u_tree.prediction_valid ;
 wire \tree_instances[11].u_tree.ready_for_next ;
 wire \tree_instances[11].u_tree.tree_state[0] ;
 wire \tree_instances[11].u_tree.tree_state[1] ;
 wire \tree_instances[11].u_tree.tree_state[2] ;
 wire \tree_instances[11].u_tree.tree_state[3] ;
 wire \tree_instances[12].u_tree.current_node_data[12] ;
 wire \tree_instances[12].u_tree.frame_id_out[0] ;
 wire \tree_instances[12].u_tree.frame_id_out[1] ;
 wire \tree_instances[12].u_tree.frame_id_out[2] ;
 wire \tree_instances[12].u_tree.frame_id_out[3] ;
 wire \tree_instances[12].u_tree.frame_id_out[4] ;
 wire \tree_instances[12].u_tree.node_data[12] ;
 wire \tree_instances[12].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[12].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[12].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[12].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[12].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[12].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[12].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[12].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[12].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[12].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[12].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[12].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[12].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[12].u_tree.pipeline_prediction[0][0] ;
 wire \tree_instances[12].u_tree.pipeline_valid[0] ;
 wire \tree_instances[12].u_tree.prediction_out ;
 wire \tree_instances[12].u_tree.prediction_valid ;
 wire \tree_instances[12].u_tree.read_enable ;
 wire \tree_instances[12].u_tree.ready_for_next ;
 wire \tree_instances[12].u_tree.tree_state[0] ;
 wire \tree_instances[12].u_tree.tree_state[1] ;
 wire \tree_instances[12].u_tree.tree_state[2] ;
 wire \tree_instances[12].u_tree.tree_state[3] ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.cache_valid ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[0] ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[1] ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[2] ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[3] ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[4] ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[5] ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[6] ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[7] ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.cached_data[12] ;
 wire \tree_instances[12].u_tree.u_tree_weight_rom.gen_tree_12.u_tree_rom.node_data[12] ;
 wire \tree_instances[13].u_tree.current_node_data[12] ;
 wire \tree_instances[13].u_tree.frame_id_out[0] ;
 wire \tree_instances[13].u_tree.frame_id_out[1] ;
 wire \tree_instances[13].u_tree.frame_id_out[2] ;
 wire \tree_instances[13].u_tree.frame_id_out[3] ;
 wire \tree_instances[13].u_tree.frame_id_out[4] ;
 wire \tree_instances[13].u_tree.node_data[12] ;
 wire \tree_instances[13].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[13].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[13].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[13].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[13].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[13].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[13].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[13].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[13].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[13].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[13].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[13].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[13].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[13].u_tree.pipeline_prediction[0][0] ;
 wire \tree_instances[13].u_tree.pipeline_valid[0] ;
 wire \tree_instances[13].u_tree.prediction_out ;
 wire \tree_instances[13].u_tree.prediction_valid ;
 wire \tree_instances[13].u_tree.read_enable ;
 wire \tree_instances[13].u_tree.ready_for_next ;
 wire \tree_instances[13].u_tree.tree_state[0] ;
 wire \tree_instances[13].u_tree.tree_state[1] ;
 wire \tree_instances[13].u_tree.tree_state[2] ;
 wire \tree_instances[13].u_tree.tree_state[3] ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.cache_valid ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[0] ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[1] ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[2] ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[3] ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[4] ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[5] ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[6] ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[7] ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.cached_data[12] ;
 wire \tree_instances[13].u_tree.u_tree_weight_rom.gen_tree_13.u_tree_rom.node_data[12] ;
 wire \tree_instances[14].u_tree.frame_id_out[0] ;
 wire \tree_instances[14].u_tree.frame_id_out[1] ;
 wire \tree_instances[14].u_tree.frame_id_out[2] ;
 wire \tree_instances[14].u_tree.frame_id_out[3] ;
 wire \tree_instances[14].u_tree.frame_id_out[4] ;
 wire \tree_instances[14].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[14].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[14].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[14].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[14].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[14].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[14].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[14].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[14].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[14].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[14].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[14].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[14].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[14].u_tree.pipeline_valid[0] ;
 wire \tree_instances[14].u_tree.prediction_valid ;
 wire \tree_instances[14].u_tree.ready_for_next ;
 wire \tree_instances[14].u_tree.tree_state[0] ;
 wire \tree_instances[14].u_tree.tree_state[1] ;
 wire \tree_instances[14].u_tree.tree_state[2] ;
 wire \tree_instances[14].u_tree.tree_state[3] ;
 wire \tree_instances[15].u_tree.frame_id_out[0] ;
 wire \tree_instances[15].u_tree.frame_id_out[1] ;
 wire \tree_instances[15].u_tree.frame_id_out[2] ;
 wire \tree_instances[15].u_tree.frame_id_out[3] ;
 wire \tree_instances[15].u_tree.frame_id_out[4] ;
 wire \tree_instances[15].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[15].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[15].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[15].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[15].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[15].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[15].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[15].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[15].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[15].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[15].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[15].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[15].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[15].u_tree.pipeline_valid[0] ;
 wire \tree_instances[15].u_tree.prediction_valid ;
 wire \tree_instances[15].u_tree.ready_for_next ;
 wire \tree_instances[15].u_tree.tree_state[0] ;
 wire \tree_instances[15].u_tree.tree_state[1] ;
 wire \tree_instances[15].u_tree.tree_state[2] ;
 wire \tree_instances[15].u_tree.tree_state[3] ;
 wire \tree_instances[16].u_tree.current_node_data[12] ;
 wire \tree_instances[16].u_tree.frame_id_out[0] ;
 wire \tree_instances[16].u_tree.frame_id_out[1] ;
 wire \tree_instances[16].u_tree.frame_id_out[2] ;
 wire \tree_instances[16].u_tree.frame_id_out[3] ;
 wire \tree_instances[16].u_tree.frame_id_out[4] ;
 wire \tree_instances[16].u_tree.node_data[12] ;
 wire \tree_instances[16].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[16].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[16].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[16].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[16].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[16].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[16].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[16].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[16].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[16].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[16].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[16].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[16].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[16].u_tree.pipeline_prediction[0][0] ;
 wire \tree_instances[16].u_tree.pipeline_valid[0] ;
 wire \tree_instances[16].u_tree.prediction_out ;
 wire \tree_instances[16].u_tree.prediction_valid ;
 wire \tree_instances[16].u_tree.read_enable ;
 wire \tree_instances[16].u_tree.ready_for_next ;
 wire \tree_instances[16].u_tree.tree_state[0] ;
 wire \tree_instances[16].u_tree.tree_state[1] ;
 wire \tree_instances[16].u_tree.tree_state[2] ;
 wire \tree_instances[16].u_tree.tree_state[3] ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.cache_valid ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[0] ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[1] ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[2] ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[3] ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[4] ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[5] ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[6] ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[7] ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.cached_data[12] ;
 wire \tree_instances[16].u_tree.u_tree_weight_rom.gen_tree_16.u_tree_rom.node_data[12] ;
 wire \tree_instances[17].u_tree.frame_id_out[0] ;
 wire \tree_instances[17].u_tree.frame_id_out[1] ;
 wire \tree_instances[17].u_tree.frame_id_out[2] ;
 wire \tree_instances[17].u_tree.frame_id_out[3] ;
 wire \tree_instances[17].u_tree.frame_id_out[4] ;
 wire \tree_instances[17].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[17].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[17].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[17].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[17].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[17].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[17].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[17].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[17].u_tree.pipeline_current_node[0][8] ;
 wire \tree_instances[17].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[17].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[17].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[17].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[17].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[17].u_tree.pipeline_valid[0] ;
 wire \tree_instances[17].u_tree.prediction_valid ;
 wire \tree_instances[17].u_tree.ready_for_next ;
 wire \tree_instances[17].u_tree.tree_state[0] ;
 wire \tree_instances[17].u_tree.tree_state[1] ;
 wire \tree_instances[17].u_tree.tree_state[2] ;
 wire \tree_instances[17].u_tree.tree_state[3] ;
 wire \tree_instances[18].u_tree.frame_id_out[0] ;
 wire \tree_instances[18].u_tree.frame_id_out[1] ;
 wire \tree_instances[18].u_tree.frame_id_out[2] ;
 wire \tree_instances[18].u_tree.frame_id_out[3] ;
 wire \tree_instances[18].u_tree.frame_id_out[4] ;
 wire \tree_instances[18].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[18].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[18].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[18].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[18].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[18].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[18].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[18].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[18].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[18].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[18].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[18].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[18].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[18].u_tree.pipeline_valid[0] ;
 wire \tree_instances[18].u_tree.prediction_valid ;
 wire \tree_instances[18].u_tree.ready_for_next ;
 wire \tree_instances[18].u_tree.tree_state[0] ;
 wire \tree_instances[18].u_tree.tree_state[1] ;
 wire \tree_instances[18].u_tree.tree_state[2] ;
 wire \tree_instances[18].u_tree.tree_state[3] ;
 wire \tree_instances[19].u_tree.frame_id_out[0] ;
 wire \tree_instances[19].u_tree.frame_id_out[1] ;
 wire \tree_instances[19].u_tree.frame_id_out[2] ;
 wire \tree_instances[19].u_tree.frame_id_out[3] ;
 wire \tree_instances[19].u_tree.frame_id_out[4] ;
 wire \tree_instances[19].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[19].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[19].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[19].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[19].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[19].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[19].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[19].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[19].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[19].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[19].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[19].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[19].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[19].u_tree.pipeline_valid[0] ;
 wire \tree_instances[19].u_tree.prediction_valid ;
 wire \tree_instances[19].u_tree.ready_for_next ;
 wire \tree_instances[19].u_tree.tree_state[0] ;
 wire \tree_instances[19].u_tree.tree_state[1] ;
 wire \tree_instances[19].u_tree.tree_state[2] ;
 wire \tree_instances[19].u_tree.tree_state[3] ;
 wire \tree_instances[1].u_tree.current_node_data[12] ;
 wire \tree_instances[1].u_tree.frame_id_out[0] ;
 wire \tree_instances[1].u_tree.frame_id_out[1] ;
 wire \tree_instances[1].u_tree.frame_id_out[2] ;
 wire \tree_instances[1].u_tree.frame_id_out[3] ;
 wire \tree_instances[1].u_tree.frame_id_out[4] ;
 wire \tree_instances[1].u_tree.node_data[12] ;
 wire \tree_instances[1].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[1].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[1].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[1].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[1].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[1].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[1].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[1].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[1].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[1].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[1].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[1].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[1].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[1].u_tree.pipeline_prediction[0][0] ;
 wire \tree_instances[1].u_tree.pipeline_valid[0] ;
 wire \tree_instances[1].u_tree.prediction_out ;
 wire \tree_instances[1].u_tree.prediction_valid ;
 wire \tree_instances[1].u_tree.read_enable ;
 wire \tree_instances[1].u_tree.ready_for_next ;
 wire \tree_instances[1].u_tree.tree_state[0] ;
 wire \tree_instances[1].u_tree.tree_state[1] ;
 wire \tree_instances[1].u_tree.tree_state[2] ;
 wire \tree_instances[1].u_tree.tree_state[3] ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.cache_valid ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[0] ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[1] ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[2] ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[3] ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[4] ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[5] ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[6] ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[7] ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.cached_data[12] ;
 wire \tree_instances[1].u_tree.u_tree_weight_rom.gen_tree_1.u_tree_rom.node_data[12] ;
 wire \tree_instances[20].u_tree.current_node_data[12] ;
 wire \tree_instances[20].u_tree.frame_id_out[0] ;
 wire \tree_instances[20].u_tree.frame_id_out[1] ;
 wire \tree_instances[20].u_tree.frame_id_out[2] ;
 wire \tree_instances[20].u_tree.frame_id_out[3] ;
 wire \tree_instances[20].u_tree.frame_id_out[4] ;
 wire \tree_instances[20].u_tree.node_data[12] ;
 wire \tree_instances[20].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[20].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[20].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[20].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[20].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[20].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[20].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[20].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[20].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[20].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[20].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[20].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[20].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[20].u_tree.pipeline_prediction[0][0] ;
 wire \tree_instances[20].u_tree.pipeline_valid[0] ;
 wire \tree_instances[20].u_tree.prediction_out ;
 wire \tree_instances[20].u_tree.prediction_valid ;
 wire \tree_instances[20].u_tree.read_enable ;
 wire \tree_instances[20].u_tree.ready_for_next ;
 wire \tree_instances[20].u_tree.tree_state[0] ;
 wire \tree_instances[20].u_tree.tree_state[1] ;
 wire \tree_instances[20].u_tree.tree_state[2] ;
 wire \tree_instances[20].u_tree.tree_state[3] ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.cache_valid ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[0] ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[1] ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[2] ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[3] ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[4] ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[5] ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[6] ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[7] ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.cached_data[12] ;
 wire \tree_instances[20].u_tree.u_tree_weight_rom.gen_tree_20.u_tree_rom.node_data[12] ;
 wire \tree_instances[2].u_tree.frame_id_out[0] ;
 wire \tree_instances[2].u_tree.frame_id_out[1] ;
 wire \tree_instances[2].u_tree.frame_id_out[2] ;
 wire \tree_instances[2].u_tree.frame_id_out[3] ;
 wire \tree_instances[2].u_tree.frame_id_out[4] ;
 wire \tree_instances[2].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[2].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[2].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[2].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[2].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[2].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[2].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[2].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[2].u_tree.pipeline_current_node[0][8] ;
 wire \tree_instances[2].u_tree.pipeline_current_node[0][9] ;
 wire \tree_instances[2].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[2].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[2].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[2].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[2].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[2].u_tree.pipeline_valid[0] ;
 wire \tree_instances[2].u_tree.prediction_valid ;
 wire \tree_instances[2].u_tree.ready_for_next ;
 wire \tree_instances[2].u_tree.tree_state[0] ;
 wire \tree_instances[2].u_tree.tree_state[1] ;
 wire \tree_instances[2].u_tree.tree_state[2] ;
 wire \tree_instances[2].u_tree.tree_state[3] ;
 wire \tree_instances[3].u_tree.current_node_data[107] ;
 wire \tree_instances[3].u_tree.frame_id_out[0] ;
 wire \tree_instances[3].u_tree.frame_id_out[1] ;
 wire \tree_instances[3].u_tree.frame_id_out[2] ;
 wire \tree_instances[3].u_tree.frame_id_out[3] ;
 wire \tree_instances[3].u_tree.frame_id_out[4] ;
 wire \tree_instances[3].u_tree.node_data[107] ;
 wire \tree_instances[3].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[3].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[3].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[3].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[3].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[3].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[3].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[3].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[3].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[3].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[3].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[3].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[3].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[3].u_tree.pipeline_prediction[0][0] ;
 wire \tree_instances[3].u_tree.pipeline_valid[0] ;
 wire \tree_instances[3].u_tree.prediction_out ;
 wire \tree_instances[3].u_tree.prediction_valid ;
 wire \tree_instances[3].u_tree.read_enable ;
 wire \tree_instances[3].u_tree.ready_for_next ;
 wire \tree_instances[3].u_tree.tree_state[0] ;
 wire \tree_instances[3].u_tree.tree_state[1] ;
 wire \tree_instances[3].u_tree.tree_state[2] ;
 wire \tree_instances[3].u_tree.tree_state[3] ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.cache_valid ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[0] ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[1] ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[2] ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[3] ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[4] ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[5] ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[6] ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[7] ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.cached_data[107] ;
 wire \tree_instances[3].u_tree.u_tree_weight_rom.gen_tree_3.u_tree_rom.node_data[107] ;
 wire \tree_instances[4].u_tree.frame_id_out[0] ;
 wire \tree_instances[4].u_tree.frame_id_out[1] ;
 wire \tree_instances[4].u_tree.frame_id_out[2] ;
 wire \tree_instances[4].u_tree.frame_id_out[3] ;
 wire \tree_instances[4].u_tree.frame_id_out[4] ;
 wire \tree_instances[4].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[4].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[4].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[4].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[4].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[4].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[4].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[4].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[4].u_tree.pipeline_current_node[0][8] ;
 wire \tree_instances[4].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[4].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[4].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[4].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[4].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[4].u_tree.pipeline_valid[0] ;
 wire \tree_instances[4].u_tree.prediction_valid ;
 wire \tree_instances[4].u_tree.ready_for_next ;
 wire \tree_instances[4].u_tree.tree_state[0] ;
 wire \tree_instances[4].u_tree.tree_state[1] ;
 wire \tree_instances[4].u_tree.tree_state[2] ;
 wire \tree_instances[4].u_tree.tree_state[3] ;
 wire \tree_instances[5].u_tree.current_node_data[107] ;
 wire \tree_instances[5].u_tree.frame_id_out[0] ;
 wire \tree_instances[5].u_tree.frame_id_out[1] ;
 wire \tree_instances[5].u_tree.frame_id_out[2] ;
 wire \tree_instances[5].u_tree.frame_id_out[3] ;
 wire \tree_instances[5].u_tree.frame_id_out[4] ;
 wire \tree_instances[5].u_tree.node_data[107] ;
 wire \tree_instances[5].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[5].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[5].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[5].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[5].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[5].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[5].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[5].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[5].u_tree.pipeline_current_node[0][8] ;
 wire \tree_instances[5].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[5].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[5].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[5].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[5].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[5].u_tree.pipeline_prediction[0][0] ;
 wire \tree_instances[5].u_tree.pipeline_valid[0] ;
 wire \tree_instances[5].u_tree.prediction_out ;
 wire \tree_instances[5].u_tree.prediction_valid ;
 wire \tree_instances[5].u_tree.read_enable ;
 wire \tree_instances[5].u_tree.ready_for_next ;
 wire \tree_instances[5].u_tree.tree_state[0] ;
 wire \tree_instances[5].u_tree.tree_state[1] ;
 wire \tree_instances[5].u_tree.tree_state[2] ;
 wire \tree_instances[5].u_tree.tree_state[3] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cache_valid ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[0] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[1] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[2] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[3] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[4] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[5] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[6] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[7] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[8] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.cached_data[107] ;
 wire \tree_instances[5].u_tree.u_tree_weight_rom.gen_tree_5.u_tree_rom.node_data[107] ;
 wire \tree_instances[6].u_tree.frame_id_out[0] ;
 wire \tree_instances[6].u_tree.frame_id_out[1] ;
 wire \tree_instances[6].u_tree.frame_id_out[2] ;
 wire \tree_instances[6].u_tree.frame_id_out[3] ;
 wire \tree_instances[6].u_tree.frame_id_out[4] ;
 wire \tree_instances[6].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[6].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[6].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[6].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[6].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[6].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[6].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[6].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[6].u_tree.pipeline_current_node[0][8] ;
 wire \tree_instances[6].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[6].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[6].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[6].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[6].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[6].u_tree.pipeline_valid[0] ;
 wire \tree_instances[6].u_tree.prediction_valid ;
 wire \tree_instances[6].u_tree.ready_for_next ;
 wire \tree_instances[6].u_tree.tree_state[0] ;
 wire \tree_instances[6].u_tree.tree_state[1] ;
 wire \tree_instances[6].u_tree.tree_state[2] ;
 wire \tree_instances[6].u_tree.tree_state[3] ;
 wire \tree_instances[7].u_tree.frame_id_out[0] ;
 wire \tree_instances[7].u_tree.frame_id_out[1] ;
 wire \tree_instances[7].u_tree.frame_id_out[2] ;
 wire \tree_instances[7].u_tree.frame_id_out[3] ;
 wire \tree_instances[7].u_tree.frame_id_out[4] ;
 wire \tree_instances[7].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[7].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[7].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[7].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[7].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[7].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[7].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[7].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[7].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[7].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[7].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[7].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[7].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[7].u_tree.pipeline_valid[0] ;
 wire \tree_instances[7].u_tree.prediction_valid ;
 wire \tree_instances[7].u_tree.ready_for_next ;
 wire \tree_instances[7].u_tree.tree_state[0] ;
 wire \tree_instances[7].u_tree.tree_state[1] ;
 wire \tree_instances[7].u_tree.tree_state[2] ;
 wire \tree_instances[7].u_tree.tree_state[3] ;
 wire \tree_instances[8].u_tree.current_node_data[12] ;
 wire \tree_instances[8].u_tree.frame_id_out[0] ;
 wire \tree_instances[8].u_tree.frame_id_out[1] ;
 wire \tree_instances[8].u_tree.frame_id_out[2] ;
 wire \tree_instances[8].u_tree.frame_id_out[3] ;
 wire \tree_instances[8].u_tree.frame_id_out[4] ;
 wire \tree_instances[8].u_tree.node_data[12] ;
 wire \tree_instances[8].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[8].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[8].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[8].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[8].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[8].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[8].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[8].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[8].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[8].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[8].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[8].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[8].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[8].u_tree.pipeline_prediction[0][0] ;
 wire \tree_instances[8].u_tree.pipeline_valid[0] ;
 wire \tree_instances[8].u_tree.prediction_out ;
 wire \tree_instances[8].u_tree.prediction_valid ;
 wire \tree_instances[8].u_tree.read_enable ;
 wire \tree_instances[8].u_tree.ready_for_next ;
 wire \tree_instances[8].u_tree.tree_state[0] ;
 wire \tree_instances[8].u_tree.tree_state[1] ;
 wire \tree_instances[8].u_tree.tree_state[2] ;
 wire \tree_instances[8].u_tree.tree_state[3] ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.cache_valid ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[0] ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[1] ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[2] ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[3] ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[4] ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[5] ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[6] ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[7] ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.cached_data[12] ;
 wire \tree_instances[8].u_tree.u_tree_weight_rom.gen_tree_8.u_tree_rom.node_data[12] ;
 wire \tree_instances[9].u_tree.frame_id_out[0] ;
 wire \tree_instances[9].u_tree.frame_id_out[1] ;
 wire \tree_instances[9].u_tree.frame_id_out[2] ;
 wire \tree_instances[9].u_tree.frame_id_out[3] ;
 wire \tree_instances[9].u_tree.frame_id_out[4] ;
 wire \tree_instances[9].u_tree.pipeline_current_node[0][0] ;
 wire \tree_instances[9].u_tree.pipeline_current_node[0][1] ;
 wire \tree_instances[9].u_tree.pipeline_current_node[0][2] ;
 wire \tree_instances[9].u_tree.pipeline_current_node[0][3] ;
 wire \tree_instances[9].u_tree.pipeline_current_node[0][4] ;
 wire \tree_instances[9].u_tree.pipeline_current_node[0][5] ;
 wire \tree_instances[9].u_tree.pipeline_current_node[0][6] ;
 wire \tree_instances[9].u_tree.pipeline_current_node[0][7] ;
 wire \tree_instances[9].u_tree.pipeline_frame_id[0][0] ;
 wire \tree_instances[9].u_tree.pipeline_frame_id[0][1] ;
 wire \tree_instances[9].u_tree.pipeline_frame_id[0][2] ;
 wire \tree_instances[9].u_tree.pipeline_frame_id[0][3] ;
 wire \tree_instances[9].u_tree.pipeline_frame_id[0][4] ;
 wire \tree_instances[9].u_tree.pipeline_valid[0] ;
 wire \tree_instances[9].u_tree.prediction_valid ;
 wire \tree_instances[9].u_tree.ready_for_next ;
 wire \tree_instances[9].u_tree.tree_state[0] ;
 wire \tree_instances[9].u_tree.tree_state[1] ;
 wire \tree_instances[9].u_tree.tree_state[2] ;
 wire \tree_instances[9].u_tree.tree_state[3] ;

 sky130_fd_sc_hd__buf_1 _3149_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][5] ),
    .X(_0705_));
 sky130_fd_sc_hd__buf_1 _3150_ (.A(_0705_),
    .X(_0706_));
 sky130_fd_sc_hd__buf_1 _3151_ (.A(_0706_),
    .X(_0707_));
 sky130_fd_sc_hd__buf_1 _3152_ (.A(_0707_),
    .X(_0708_));
 sky130_fd_sc_hd__buf_1 _3153_ (.A(_0708_),
    .X(_0709_));
 sky130_fd_sc_hd__buf_1 _3154_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][2] ),
    .X(_0710_));
 sky130_fd_sc_hd__buf_1 _3155_ (.A(_0710_),
    .X(_0711_));
 sky130_fd_sc_hd__buf_1 _3156_ (.A(_0711_),
    .X(_0712_));
 sky130_fd_sc_hd__buf_1 _3157_ (.A(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__buf_1 _3158_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][4] ),
    .X(_0714_));
 sky130_fd_sc_hd__buf_1 _3159_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][3] ),
    .X(_0715_));
 sky130_fd_sc_hd__buf_1 _3160_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][1] ),
    .X(_0716_));
 sky130_fd_sc_hd__buf_1 _3161_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][0] ),
    .X(_0717_));
 sky130_fd_sc_hd__or3_2 _3162_ (.A(_0715_),
    .B(_0716_),
    .C(_0717_),
    .X(_0718_));
 sky130_fd_sc_hd__or2_2 _3163_ (.A(_0714_),
    .B(_0718_),
    .X(_0719_));
 sky130_fd_sc_hd__or2_2 _3164_ (.A(_0713_),
    .B(_0719_),
    .X(_0720_));
 sky130_fd_sc_hd__buf_1 _3165_ (.A(_0720_),
    .X(_0721_));
 sky130_fd_sc_hd__inv_2 _3166_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][8] ),
    .Y(_0722_));
 sky130_fd_sc_hd__buf_1 _3167_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][6] ),
    .X(_0723_));
 sky130_fd_sc_hd__buf_1 _3168_ (.A(_0723_),
    .X(_0724_));
 sky130_fd_sc_hd__buf_1 _3169_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][7] ),
    .X(_0725_));
 sky130_fd_sc_hd__buf_1 _3170_ (.A(_0725_),
    .X(_0726_));
 sky130_fd_sc_hd__nor2_2 _3171_ (.A(_0724_),
    .B(_0726_),
    .Y(_0727_));
 sky130_fd_sc_hd__nand2_2 _3172_ (.A(_0722_),
    .B(_0727_),
    .Y(_0728_));
 sky130_fd_sc_hd__buf_1 _3173_ (.A(\tree_instances[4].u_tree.tree_state[2] ),
    .X(_0729_));
 sky130_fd_sc_hd__o31a_2 _3174_ (.A1(_0709_),
    .A2(_0721_),
    .A3(_0728_),
    .B1(_0729_),
    .X(_0033_));
 sky130_fd_sc_hd__inv_2 _3175_ (.A(feature_valid),
    .Y(_0730_));
 sky130_fd_sc_hd__buf_1 _3176_ (.A(_0730_),
    .X(_0731_));
 sky130_fd_sc_hd__buf_1 _3177_ (.A(_0731_),
    .X(_0732_));
 sky130_fd_sc_hd__buf_1 _3178_ (.A(_0732_),
    .X(_0733_));
 sky130_fd_sc_hd__or2_2 _3179_ (.A(_0733_),
    .B(\tree_instances[14].u_tree.pipeline_valid[0] ),
    .X(_0734_));
 sky130_fd_sc_hd__buf_1 _3180_ (.A(\tree_instances[14].u_tree.tree_state[3] ),
    .X(_0735_));
 sky130_fd_sc_hd__a21o_2 _3181_ (.A1(\tree_instances[14].u_tree.tree_state[0] ),
    .A2(_0734_),
    .B1(_0735_),
    .X(_0055_));
 sky130_fd_sc_hd__or2_2 _3182_ (.A(_0733_),
    .B(\tree_instances[0].u_tree.pipeline_valid[0] ),
    .X(_0736_));
 sky130_fd_sc_hd__buf_1 _3183_ (.A(\tree_instances[0].u_tree.tree_state[3] ),
    .X(_0737_));
 sky130_fd_sc_hd__a21o_2 _3184_ (.A1(\tree_instances[0].u_tree.tree_state[0] ),
    .A2(_0736_),
    .B1(_0737_),
    .X(_0045_));
 sky130_fd_sc_hd__buf_1 _3185_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][2] ),
    .X(_0738_));
 sky130_fd_sc_hd__or2_2 _3186_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][3] ),
    .B(_0738_),
    .X(_0739_));
 sky130_fd_sc_hd__or2_2 _3187_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][1] ),
    .B(\tree_instances[18].u_tree.pipeline_current_node[0][0] ),
    .X(_0740_));
 sky130_fd_sc_hd__buf_1 _3188_ (.A(_0740_),
    .X(_0741_));
 sky130_fd_sc_hd__or2_2 _3189_ (.A(_0739_),
    .B(_0741_),
    .X(_0742_));
 sky130_fd_sc_hd__buf_1 _3190_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][7] ),
    .X(_0743_));
 sky130_fd_sc_hd__or2_2 _3191_ (.A(_0743_),
    .B(\tree_instances[18].u_tree.pipeline_current_node[0][6] ),
    .X(_0744_));
 sky130_fd_sc_hd__buf_1 _3192_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][5] ),
    .X(_0745_));
 sky130_fd_sc_hd__buf_1 _3193_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][4] ),
    .X(_0746_));
 sky130_fd_sc_hd__buf_1 _3194_ (.A(_0746_),
    .X(_0747_));
 sky130_fd_sc_hd__or2_2 _3195_ (.A(_0745_),
    .B(_0747_),
    .X(_0748_));
 sky130_fd_sc_hd__buf_1 _3196_ (.A(_0748_),
    .X(_0749_));
 sky130_fd_sc_hd__buf_1 _3197_ (.A(_0749_),
    .X(_0750_));
 sky130_fd_sc_hd__buf_1 _3198_ (.A(\tree_instances[18].u_tree.tree_state[2] ),
    .X(_0751_));
 sky130_fd_sc_hd__o31a_2 _3199_ (.A1(_0742_),
    .A2(_0744_),
    .A3(_0750_),
    .B1(_0751_),
    .X(_0021_));
 sky130_fd_sc_hd__or2_2 _3200_ (.A(_0733_),
    .B(\tree_instances[18].u_tree.pipeline_valid[0] ),
    .X(_0752_));
 sky130_fd_sc_hd__buf_1 _3201_ (.A(\tree_instances[18].u_tree.tree_state[3] ),
    .X(_0753_));
 sky130_fd_sc_hd__a21o_2 _3202_ (.A1(\tree_instances[18].u_tree.tree_state[0] ),
    .A2(_0752_),
    .B1(_0753_),
    .X(_0063_));
 sky130_fd_sc_hd__or2_2 _3203_ (.A(_0733_),
    .B(\tree_instances[2].u_tree.pipeline_valid[0] ),
    .X(_0754_));
 sky130_fd_sc_hd__buf_1 _3204_ (.A(\tree_instances[2].u_tree.tree_state[3] ),
    .X(_0755_));
 sky130_fd_sc_hd__a21o_2 _3205_ (.A1(\tree_instances[2].u_tree.tree_state[0] ),
    .A2(_0754_),
    .B1(_0755_),
    .X(_0071_));
 sky130_fd_sc_hd__buf_1 _3206_ (.A(\tree_instances[20].u_tree.tree_state[2] ),
    .X(_0756_));
 sky130_fd_sc_hd__buf_1 _3207_ (.A(_0756_),
    .X(_0757_));
 sky130_fd_sc_hd__buf_1 _3208_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][6] ),
    .X(_0758_));
 sky130_fd_sc_hd__nor2_2 _3209_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][7] ),
    .B(_0758_),
    .Y(_0759_));
 sky130_fd_sc_hd__buf_1 _3210_ (.A(_0759_),
    .X(_0760_));
 sky130_fd_sc_hd__buf_1 _3211_ (.A(_0760_),
    .X(_0761_));
 sky130_fd_sc_hd__or2_2 _3212_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][1] ),
    .B(\tree_instances[20].u_tree.pipeline_current_node[0][0] ),
    .X(_0762_));
 sky130_fd_sc_hd__buf_1 _3213_ (.A(_0762_),
    .X(_0763_));
 sky130_fd_sc_hd__buf_1 _3214_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][3] ),
    .X(_0764_));
 sky130_fd_sc_hd__buf_1 _3215_ (.A(_0764_),
    .X(_0765_));
 sky130_fd_sc_hd__buf_1 _3216_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][2] ),
    .X(_0766_));
 sky130_fd_sc_hd__buf_1 _3217_ (.A(_0766_),
    .X(_0767_));
 sky130_fd_sc_hd__or2_2 _3218_ (.A(_0765_),
    .B(_0767_),
    .X(_0768_));
 sky130_fd_sc_hd__buf_1 _3219_ (.A(_0768_),
    .X(_0769_));
 sky130_fd_sc_hd__nor2_2 _3220_ (.A(_0763_),
    .B(_0769_),
    .Y(_0770_));
 sky130_fd_sc_hd__nor2_2 _3221_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][5] ),
    .B(\tree_instances[20].u_tree.pipeline_current_node[0][4] ),
    .Y(_0771_));
 sky130_fd_sc_hd__buf_1 _3222_ (.A(_0771_),
    .X(_0772_));
 sky130_fd_sc_hd__buf_1 _3223_ (.A(_0772_),
    .X(_0773_));
 sky130_fd_sc_hd__buf_1 _3224_ (.A(_0773_),
    .X(_0774_));
 sky130_fd_sc_hd__a41o_2 _3225_ (.A1(_0757_),
    .A2(_0761_),
    .A3(_0770_),
    .A4(_0774_),
    .B1(\tree_instances[20].u_tree.tree_state[1] ),
    .X(_0070_));
 sky130_fd_sc_hd__buf_1 _3226_ (.A(\tree_instances[17].u_tree.tree_state[2] ),
    .X(_0775_));
 sky130_fd_sc_hd__buf_1 _3227_ (.A(_0775_),
    .X(_0776_));
 sky130_fd_sc_hd__nor2_2 _3228_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][8] ),
    .B(\tree_instances[17].u_tree.pipeline_current_node[0][7] ),
    .Y(_0777_));
 sky130_fd_sc_hd__buf_1 _3229_ (.A(_0777_),
    .X(_0778_));
 sky130_fd_sc_hd__buf_1 _3230_ (.A(_0778_),
    .X(_0779_));
 sky130_fd_sc_hd__buf_1 _3231_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][2] ),
    .X(_0780_));
 sky130_fd_sc_hd__buf_1 _3232_ (.A(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__buf_1 _3233_ (.A(_0781_),
    .X(_0782_));
 sky130_fd_sc_hd__inv_2 _3234_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][3] ),
    .Y(_0783_));
 sky130_fd_sc_hd__buf_1 _3235_ (.A(_0783_),
    .X(_0784_));
 sky130_fd_sc_hd__buf_1 _3236_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][1] ),
    .X(_0785_));
 sky130_fd_sc_hd__buf_1 _3237_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][0] ),
    .X(_0786_));
 sky130_fd_sc_hd__nor2_2 _3238_ (.A(_0785_),
    .B(_0786_),
    .Y(_0787_));
 sky130_fd_sc_hd__nand2_2 _3239_ (.A(_0784_),
    .B(_0787_),
    .Y(_0788_));
 sky130_fd_sc_hd__or2_2 _3240_ (.A(_0782_),
    .B(_0788_),
    .X(_0789_));
 sky130_fd_sc_hd__inv_2 _3241_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][6] ),
    .Y(_0790_));
 sky130_fd_sc_hd__buf_1 _3242_ (.A(_0790_),
    .X(_0791_));
 sky130_fd_sc_hd__buf_1 _3243_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][5] ),
    .X(_0792_));
 sky130_fd_sc_hd__buf_1 _3244_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][4] ),
    .X(_0793_));
 sky130_fd_sc_hd__buf_1 _3245_ (.A(_0793_),
    .X(_0794_));
 sky130_fd_sc_hd__nor2_2 _3246_ (.A(_0792_),
    .B(_0794_),
    .Y(_0795_));
 sky130_fd_sc_hd__buf_1 _3247_ (.A(_0795_),
    .X(_0796_));
 sky130_fd_sc_hd__nand2_2 _3248_ (.A(_0791_),
    .B(_0796_),
    .Y(_0797_));
 sky130_fd_sc_hd__nor2_2 _3249_ (.A(_0789_),
    .B(_0797_),
    .Y(_0798_));
 sky130_fd_sc_hd__a31o_2 _3250_ (.A1(_0776_),
    .A2(_0779_),
    .A3(_0798_),
    .B1(\tree_instances[17].u_tree.tree_state[1] ),
    .X(_0062_));
 sky130_fd_sc_hd__buf_1 _3251_ (.A(\tree_instances[3].u_tree.tree_state[3] ),
    .X(_0799_));
 sky130_fd_sc_hd__o21ai_2 _3252_ (.A1(_0732_),
    .A2(\tree_instances[3].u_tree.pipeline_valid[0] ),
    .B1(\tree_instances[3].u_tree.tree_state[0] ),
    .Y(_0800_));
 sky130_fd_sc_hd__or2b_2 _3253_ (.A(_0799_),
    .B_N(_0800_),
    .X(_0801_));
 sky130_fd_sc_hd__buf_1 _3254_ (.A(_0801_),
    .X(_0073_));
 sky130_fd_sc_hd__buf_1 _3255_ (.A(\tree_instances[2].u_tree.tree_state[2] ),
    .X(_0802_));
 sky130_fd_sc_hd__inv_2 _3256_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][3] ),
    .Y(_0803_));
 sky130_fd_sc_hd__nand2_2 _3257_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][6] ),
    .B(\tree_instances[2].u_tree.pipeline_current_node[0][7] ),
    .Y(_0804_));
 sky130_fd_sc_hd__nand2_2 _3258_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][5] ),
    .B(\tree_instances[2].u_tree.pipeline_current_node[0][4] ),
    .Y(_0805_));
 sky130_fd_sc_hd__or2_2 _3259_ (.A(_0804_),
    .B(_0805_),
    .X(_0806_));
 sky130_fd_sc_hd__inv_2 _3260_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][8] ),
    .Y(_0807_));
 sky130_fd_sc_hd__inv_2 _3261_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][9] ),
    .Y(_0808_));
 sky130_fd_sc_hd__o211a_2 _3262_ (.A1(_0803_),
    .A2(_0806_),
    .B1(_0807_),
    .C1(_0808_),
    .X(_0809_));
 sky130_fd_sc_hd__buf_1 _3263_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][5] ),
    .X(_0810_));
 sky130_fd_sc_hd__buf_1 _3264_ (.A(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__buf_1 _3265_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][4] ),
    .X(_0812_));
 sky130_fd_sc_hd__buf_1 _3266_ (.A(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__buf_1 _3267_ (.A(_0813_),
    .X(_0814_));
 sky130_fd_sc_hd__nor2_2 _3268_ (.A(_0811_),
    .B(_0814_),
    .Y(_0815_));
 sky130_fd_sc_hd__buf_1 _3269_ (.A(_0815_),
    .X(_0816_));
 sky130_fd_sc_hd__buf_1 _3270_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][6] ),
    .X(_0817_));
 sky130_fd_sc_hd__buf_1 _3271_ (.A(_0817_),
    .X(_0818_));
 sky130_fd_sc_hd__nor2_2 _3272_ (.A(_0818_),
    .B(\tree_instances[2].u_tree.pipeline_current_node[0][7] ),
    .Y(_0819_));
 sky130_fd_sc_hd__nand2_2 _3273_ (.A(_0816_),
    .B(_0819_),
    .Y(_0820_));
 sky130_fd_sc_hd__buf_1 _3274_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][2] ),
    .X(_0821_));
 sky130_fd_sc_hd__or2_2 _3275_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][1] ),
    .B(_0821_),
    .X(_0822_));
 sky130_fd_sc_hd__buf_1 _3276_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][0] ),
    .X(_0823_));
 sky130_fd_sc_hd__buf_1 _3277_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][3] ),
    .X(_0824_));
 sky130_fd_sc_hd__buf_1 _3278_ (.A(_0824_),
    .X(_0825_));
 sky130_fd_sc_hd__or2_2 _3279_ (.A(_0823_),
    .B(_0825_),
    .X(_0826_));
 sky130_fd_sc_hd__or2_2 _3280_ (.A(_0822_),
    .B(_0826_),
    .X(_0827_));
 sky130_fd_sc_hd__nor2_2 _3281_ (.A(_0820_),
    .B(_0827_),
    .Y(_0828_));
 sky130_fd_sc_hd__a31o_2 _3282_ (.A1(_0802_),
    .A2(_0809_),
    .A3(_0828_),
    .B1(\tree_instances[2].u_tree.tree_state[1] ),
    .X(_0072_));
 sky130_fd_sc_hd__buf_1 _3283_ (.A(\tree_instances[12].u_tree.tree_state[3] ),
    .X(_0829_));
 sky130_fd_sc_hd__o21ai_2 _3284_ (.A1(_0731_),
    .A2(\tree_instances[12].u_tree.pipeline_valid[0] ),
    .B1(\tree_instances[12].u_tree.tree_state[0] ),
    .Y(_0830_));
 sky130_fd_sc_hd__or2b_2 _3285_ (.A(_0829_),
    .B_N(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__buf_1 _3286_ (.A(_0831_),
    .X(_0051_));
 sky130_fd_sc_hd__or2_2 _3287_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][5] ),
    .B(\tree_instances[12].u_tree.pipeline_current_node[0][4] ),
    .X(_0832_));
 sky130_fd_sc_hd__buf_1 _3288_ (.A(_0832_),
    .X(_0833_));
 sky130_fd_sc_hd__buf_1 _3289_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][0] ),
    .X(_0834_));
 sky130_fd_sc_hd__nor2_2 _3290_ (.A(_0834_),
    .B(\tree_instances[12].u_tree.pipeline_current_node[0][3] ),
    .Y(_0835_));
 sky130_fd_sc_hd__buf_1 _3291_ (.A(_0835_),
    .X(_0836_));
 sky130_fd_sc_hd__buf_1 _3292_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][1] ),
    .X(_0837_));
 sky130_fd_sc_hd__buf_1 _3293_ (.A(_0837_),
    .X(_0838_));
 sky130_fd_sc_hd__buf_1 _3294_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][2] ),
    .X(_0839_));
 sky130_fd_sc_hd__buf_1 _3295_ (.A(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__nor2_2 _3296_ (.A(_0838_),
    .B(_0840_),
    .Y(_0841_));
 sky130_fd_sc_hd__nand2_2 _3297_ (.A(_0836_),
    .B(_0841_),
    .Y(_0842_));
 sky130_fd_sc_hd__buf_1 _3298_ (.A(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__or2_2 _3299_ (.A(_0833_),
    .B(_0843_),
    .X(_0844_));
 sky130_fd_sc_hd__buf_1 _3300_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][6] ),
    .X(_0845_));
 sky130_fd_sc_hd__buf_1 _3301_ (.A(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__or2_2 _3302_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][7] ),
    .B(_0846_),
    .X(_0847_));
 sky130_fd_sc_hd__o21a_2 _3303_ (.A1(_0844_),
    .A2(_0847_),
    .B1(\tree_instances[12].u_tree.tree_state[2] ),
    .X(_0009_));
 sky130_fd_sc_hd__or2_2 _3304_ (.A(_0733_),
    .B(\tree_instances[4].u_tree.pipeline_valid[0] ),
    .X(_0848_));
 sky130_fd_sc_hd__buf_1 _3305_ (.A(\tree_instances[4].u_tree.tree_state[3] ),
    .X(_0849_));
 sky130_fd_sc_hd__a21o_2 _3306_ (.A1(\tree_instances[4].u_tree.tree_state[0] ),
    .A2(_0848_),
    .B1(_0849_),
    .X(_0075_));
 sky130_fd_sc_hd__buf_1 _3307_ (.A(\tree_instances[3].u_tree.tree_state[2] ),
    .X(_0850_));
 sky130_fd_sc_hd__buf_1 _3308_ (.A(_0850_),
    .X(_0851_));
 sky130_fd_sc_hd__buf_1 _3309_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][4] ),
    .X(_0852_));
 sky130_fd_sc_hd__nor2_2 _3310_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][5] ),
    .B(_0852_),
    .Y(_0853_));
 sky130_fd_sc_hd__buf_1 _3311_ (.A(_0853_),
    .X(_0854_));
 sky130_fd_sc_hd__buf_1 _3312_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][1] ),
    .X(_0855_));
 sky130_fd_sc_hd__or2_2 _3313_ (.A(_0855_),
    .B(\tree_instances[3].u_tree.pipeline_current_node[0][3] ),
    .X(_0856_));
 sky130_fd_sc_hd__buf_1 _3314_ (.A(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__buf_1 _3315_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][2] ),
    .X(_0858_));
 sky130_fd_sc_hd__or2_2 _3316_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][0] ),
    .B(_0858_),
    .X(_0859_));
 sky130_fd_sc_hd__buf_1 _3317_ (.A(_0859_),
    .X(_0860_));
 sky130_fd_sc_hd__nor2_2 _3318_ (.A(_0857_),
    .B(_0860_),
    .Y(_0861_));
 sky130_fd_sc_hd__buf_1 _3319_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][6] ),
    .X(_0862_));
 sky130_fd_sc_hd__nor2_2 _3320_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][7] ),
    .B(_0862_),
    .Y(_0863_));
 sky130_fd_sc_hd__buf_1 _3321_ (.A(_0863_),
    .X(_0864_));
 sky130_fd_sc_hd__a41o_2 _3322_ (.A1(_0851_),
    .A2(_0854_),
    .A3(_0861_),
    .A4(_0864_),
    .B1(\tree_instances[3].u_tree.tree_state[1] ),
    .X(_0074_));
 sky130_fd_sc_hd__buf_1 _3323_ (.A(\tree_instances[1].u_tree.tree_state[2] ),
    .X(_0865_));
 sky130_fd_sc_hd__buf_1 _3324_ (.A(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__buf_1 _3325_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][1] ),
    .X(_0867_));
 sky130_fd_sc_hd__buf_1 _3326_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][3] ),
    .X(_0868_));
 sky130_fd_sc_hd__or2_2 _3327_ (.A(_0867_),
    .B(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__buf_1 _3328_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][0] ),
    .X(_0870_));
 sky130_fd_sc_hd__buf_1 _3329_ (.A(_0870_),
    .X(_0871_));
 sky130_fd_sc_hd__buf_1 _3330_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][2] ),
    .X(_0872_));
 sky130_fd_sc_hd__or2_2 _3331_ (.A(_0871_),
    .B(_0872_),
    .X(_0873_));
 sky130_fd_sc_hd__or2_2 _3332_ (.A(_0869_),
    .B(_0873_),
    .X(_0874_));
 sky130_fd_sc_hd__buf_1 _3333_ (.A(_0874_),
    .X(_0875_));
 sky130_fd_sc_hd__buf_1 _3334_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][7] ),
    .X(_0876_));
 sky130_fd_sc_hd__buf_1 _3335_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][4] ),
    .X(_0877_));
 sky130_fd_sc_hd__buf_1 _3336_ (.A(_0877_),
    .X(_0878_));
 sky130_fd_sc_hd__buf_1 _3337_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][5] ),
    .X(_0879_));
 sky130_fd_sc_hd__or2_2 _3338_ (.A(_0878_),
    .B(_0879_),
    .X(_0880_));
 sky130_fd_sc_hd__buf_1 _3339_ (.A(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__or3_2 _3340_ (.A(_0876_),
    .B(\tree_instances[1].u_tree.pipeline_current_node[0][6] ),
    .C(_0881_),
    .X(_0882_));
 sky130_fd_sc_hd__nor2_2 _3341_ (.A(_0875_),
    .B(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__a21o_2 _3342_ (.A1(_0866_),
    .A2(_0883_),
    .B1(\tree_instances[1].u_tree.tree_state[1] ),
    .X(_0068_));
 sky130_fd_sc_hd__buf_1 _3343_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][3] ),
    .X(_0884_));
 sky130_fd_sc_hd__buf_1 _3344_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][4] ),
    .X(_0885_));
 sky130_fd_sc_hd__or2_2 _3345_ (.A(_0884_),
    .B(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__buf_1 _3346_ (.A(_0886_),
    .X(_0887_));
 sky130_fd_sc_hd__inv_2 _3347_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][0] ),
    .Y(_0888_));
 sky130_fd_sc_hd__buf_1 _3348_ (.A(_0888_),
    .X(_0889_));
 sky130_fd_sc_hd__buf_1 _3349_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][1] ),
    .X(_0890_));
 sky130_fd_sc_hd__buf_1 _3350_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][2] ),
    .X(_0891_));
 sky130_fd_sc_hd__nor2_2 _3351_ (.A(_0890_),
    .B(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__nand2_2 _3352_ (.A(_0889_),
    .B(_0892_),
    .Y(_0893_));
 sky130_fd_sc_hd__nor2_2 _3353_ (.A(_0887_),
    .B(_0893_),
    .Y(_0894_));
 sky130_fd_sc_hd__inv_2 _3354_ (.A(_0894_),
    .Y(_0895_));
 sky130_fd_sc_hd__inv_2 _3355_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][7] ),
    .Y(_0896_));
 sky130_fd_sc_hd__buf_1 _3356_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][5] ),
    .X(_0897_));
 sky130_fd_sc_hd__buf_1 _3357_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][6] ),
    .X(_0898_));
 sky130_fd_sc_hd__nor2_2 _3358_ (.A(_0897_),
    .B(_0898_),
    .Y(_0899_));
 sky130_fd_sc_hd__nand2_2 _3359_ (.A(_0896_),
    .B(_0899_),
    .Y(_0900_));
 sky130_fd_sc_hd__buf_1 _3360_ (.A(\tree_instances[19].u_tree.tree_state[2] ),
    .X(_0901_));
 sky130_fd_sc_hd__o21a_2 _3361_ (.A1(_0895_),
    .A2(_0900_),
    .B1(_0901_),
    .X(_0023_));
 sky130_fd_sc_hd__or2_2 _3362_ (.A(_0732_),
    .B(\tree_instances[5].u_tree.pipeline_valid[0] ),
    .X(_0902_));
 sky130_fd_sc_hd__buf_1 _3363_ (.A(\tree_instances[5].u_tree.tree_state[3] ),
    .X(_0903_));
 sky130_fd_sc_hd__a21o_2 _3364_ (.A1(\tree_instances[5].u_tree.tree_state[0] ),
    .A2(_0902_),
    .B1(_0903_),
    .X(_0077_));
 sky130_fd_sc_hd__inv_2 _3365_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][5] ),
    .Y(_0904_));
 sky130_fd_sc_hd__buf_1 _3366_ (.A(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__buf_1 _3367_ (.A(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__buf_1 _3368_ (.A(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__nor2_2 _3369_ (.A(_0721_),
    .B(_0728_),
    .Y(_0908_));
 sky130_fd_sc_hd__a31o_2 _3370_ (.A1(_0907_),
    .A2(_0729_),
    .A3(_0908_),
    .B1(\tree_instances[4].u_tree.tree_state[1] ),
    .X(_0076_));
 sky130_fd_sc_hd__buf_1 _3371_ (.A(\tree_instances[17].u_tree.tree_state[3] ),
    .X(_0909_));
 sky130_fd_sc_hd__o21a_2 _3372_ (.A1(_0732_),
    .A2(\tree_instances[17].u_tree.pipeline_valid[0] ),
    .B1(\tree_instances[17].u_tree.tree_state[0] ),
    .X(_0910_));
 sky130_fd_sc_hd__or2_2 _3373_ (.A(_0909_),
    .B(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__buf_1 _3374_ (.A(_0911_),
    .X(_0061_));
 sky130_fd_sc_hd__buf_1 _3375_ (.A(\tree_instances[16].u_tree.tree_state[2] ),
    .X(_0912_));
 sky130_fd_sc_hd__buf_1 _3376_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][7] ),
    .X(_0913_));
 sky130_fd_sc_hd__buf_1 _3377_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][6] ),
    .X(_0914_));
 sky130_fd_sc_hd__buf_1 _3378_ (.A(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__nor2_2 _3379_ (.A(_0913_),
    .B(_0915_),
    .Y(_0916_));
 sky130_fd_sc_hd__buf_1 _3380_ (.A(_0916_),
    .X(_0917_));
 sky130_fd_sc_hd__buf_1 _3381_ (.A(_0917_),
    .X(_0918_));
 sky130_fd_sc_hd__or2_2 _3382_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][1] ),
    .B(\tree_instances[16].u_tree.pipeline_current_node[0][0] ),
    .X(_0919_));
 sky130_fd_sc_hd__buf_1 _3383_ (.A(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__or2_2 _3384_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][3] ),
    .B(\tree_instances[16].u_tree.pipeline_current_node[0][2] ),
    .X(_0921_));
 sky130_fd_sc_hd__buf_1 _3385_ (.A(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__nor2_2 _3386_ (.A(_0920_),
    .B(_0922_),
    .Y(_0923_));
 sky130_fd_sc_hd__buf_1 _3387_ (.A(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__buf_1 _3388_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][5] ),
    .X(_0925_));
 sky130_fd_sc_hd__buf_1 _3389_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][4] ),
    .X(_0926_));
 sky130_fd_sc_hd__buf_1 _3390_ (.A(_0926_),
    .X(_0927_));
 sky130_fd_sc_hd__nor2_2 _3391_ (.A(_0925_),
    .B(_0927_),
    .Y(_0928_));
 sky130_fd_sc_hd__buf_1 _3392_ (.A(_0928_),
    .X(_0929_));
 sky130_fd_sc_hd__buf_1 _3393_ (.A(_0929_),
    .X(_0930_));
 sky130_fd_sc_hd__a41o_2 _3394_ (.A1(_0912_),
    .A2(_0918_),
    .A3(_0924_),
    .A4(_0930_),
    .B1(\tree_instances[16].u_tree.tree_state[1] ),
    .X(_0060_));
 sky130_fd_sc_hd__or2_2 _3395_ (.A(_0732_),
    .B(\tree_instances[6].u_tree.pipeline_valid[0] ),
    .X(_0931_));
 sky130_fd_sc_hd__buf_1 _3396_ (.A(\tree_instances[6].u_tree.tree_state[3] ),
    .X(_0932_));
 sky130_fd_sc_hd__a21o_2 _3397_ (.A1(\tree_instances[6].u_tree.tree_state[0] ),
    .A2(_0931_),
    .B1(_0932_),
    .X(_0079_));
 sky130_fd_sc_hd__buf_1 _3398_ (.A(\tree_instances[5].u_tree.tree_state[2] ),
    .X(_0933_));
 sky130_fd_sc_hd__buf_1 _3399_ (.A(_0933_),
    .X(_0934_));
 sky130_fd_sc_hd__or2_2 _3400_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][0] ),
    .B(\tree_instances[5].u_tree.pipeline_current_node[0][1] ),
    .X(_0935_));
 sky130_fd_sc_hd__buf_1 _3401_ (.A(_0935_),
    .X(_0936_));
 sky130_fd_sc_hd__buf_1 _3402_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][3] ),
    .X(_0937_));
 sky130_fd_sc_hd__buf_1 _3403_ (.A(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__buf_1 _3404_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][2] ),
    .X(_0939_));
 sky130_fd_sc_hd__buf_1 _3405_ (.A(_0939_),
    .X(_0940_));
 sky130_fd_sc_hd__or2_2 _3406_ (.A(_0938_),
    .B(_0940_),
    .X(_0941_));
 sky130_fd_sc_hd__buf_1 _3407_ (.A(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__nor2_2 _3408_ (.A(_0936_),
    .B(_0942_),
    .Y(_0943_));
 sky130_fd_sc_hd__buf_1 _3409_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][7] ),
    .X(_0944_));
 sky130_fd_sc_hd__buf_1 _3410_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][8] ),
    .X(_0945_));
 sky130_fd_sc_hd__nor2_2 _3411_ (.A(_0944_),
    .B(_0945_),
    .Y(_0946_));
 sky130_fd_sc_hd__buf_1 _3412_ (.A(_0946_),
    .X(_0947_));
 sky130_fd_sc_hd__or2_2 _3413_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][4] ),
    .B(\tree_instances[5].u_tree.pipeline_current_node[0][5] ),
    .X(_0948_));
 sky130_fd_sc_hd__buf_1 _3414_ (.A(_0948_),
    .X(_0949_));
 sky130_fd_sc_hd__nor2_2 _3415_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][6] ),
    .B(_0949_),
    .Y(_0950_));
 sky130_fd_sc_hd__a41o_2 _3416_ (.A1(_0934_),
    .A2(_0943_),
    .A3(_0947_),
    .A4(_0950_),
    .B1(\tree_instances[5].u_tree.tree_state[1] ),
    .X(_0078_));
 sky130_fd_sc_hd__inv_2 _3417_ (.A(\tree_instances[11].u_tree.tree_state[3] ),
    .Y(_0951_));
 sky130_fd_sc_hd__o21ai_2 _3418_ (.A1(_0733_),
    .A2(\tree_instances[11].u_tree.pipeline_valid[0] ),
    .B1(\tree_instances[11].u_tree.tree_state[0] ),
    .Y(_0952_));
 sky130_fd_sc_hd__nand2_2 _3419_ (.A(_0951_),
    .B(_0952_),
    .Y(_0049_));
 sky130_fd_sc_hd__inv_2 _3420_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][7] ),
    .Y(_0953_));
 sky130_fd_sc_hd__nor2_2 _3421_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][5] ),
    .B(\tree_instances[13].u_tree.pipeline_current_node[0][6] ),
    .Y(_0954_));
 sky130_fd_sc_hd__nand2_2 _3422_ (.A(_0953_),
    .B(_0954_),
    .Y(_0955_));
 sky130_fd_sc_hd__buf_1 _3423_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][2] ),
    .X(_0956_));
 sky130_fd_sc_hd__buf_1 _3424_ (.A(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__buf_1 _3425_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][1] ),
    .X(_0958_));
 sky130_fd_sc_hd__or3_2 _3426_ (.A(_0958_),
    .B(\tree_instances[13].u_tree.pipeline_current_node[0][0] ),
    .C(\tree_instances[13].u_tree.pipeline_current_node[0][3] ),
    .X(_0959_));
 sky130_fd_sc_hd__buf_1 _3427_ (.A(_0959_),
    .X(_0960_));
 sky130_fd_sc_hd__nor2_2 _3428_ (.A(_0957_),
    .B(_0960_),
    .Y(_0961_));
 sky130_fd_sc_hd__inv_2 _3429_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][4] ),
    .Y(_0962_));
 sky130_fd_sc_hd__buf_1 _3430_ (.A(_0962_),
    .X(_0963_));
 sky130_fd_sc_hd__buf_1 _3431_ (.A(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__and3b_2 _3432_ (.A_N(_0955_),
    .B(_0961_),
    .C(_0964_),
    .X(_0965_));
 sky130_fd_sc_hd__and2b_2 _3433_ (.A_N(_0965_),
    .B(\tree_instances[13].u_tree.tree_state[2] ),
    .X(_0966_));
 sky130_fd_sc_hd__buf_1 _3434_ (.A(_0966_),
    .X(_0011_));
 sky130_fd_sc_hd__buf_1 _3435_ (.A(\tree_instances[13].u_tree.tree_state[2] ),
    .X(_0967_));
 sky130_fd_sc_hd__buf_1 _3436_ (.A(_0967_),
    .X(_0968_));
 sky130_fd_sc_hd__a21o_2 _3437_ (.A1(_0968_),
    .A2(_0965_),
    .B1(\tree_instances[13].u_tree.tree_state[1] ),
    .X(_0054_));
 sky130_fd_sc_hd__or2_2 _3438_ (.A(_0733_),
    .B(\tree_instances[7].u_tree.pipeline_valid[0] ),
    .X(_0969_));
 sky130_fd_sc_hd__buf_1 _3439_ (.A(\tree_instances[7].u_tree.tree_state[3] ),
    .X(_0970_));
 sky130_fd_sc_hd__a21o_2 _3440_ (.A1(\tree_instances[7].u_tree.tree_state[0] ),
    .A2(_0969_),
    .B1(_0970_),
    .X(_0081_));
 sky130_fd_sc_hd__buf_1 _3441_ (.A(\tree_instances[6].u_tree.tree_state[2] ),
    .X(_0971_));
 sky130_fd_sc_hd__buf_1 _3442_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][5] ),
    .X(_0972_));
 sky130_fd_sc_hd__buf_1 _3443_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][4] ),
    .X(_0973_));
 sky130_fd_sc_hd__buf_1 _3444_ (.A(_0973_),
    .X(_0974_));
 sky130_fd_sc_hd__or2_2 _3445_ (.A(_0972_),
    .B(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__buf_1 _3446_ (.A(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__buf_1 _3447_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][1] ),
    .X(_0977_));
 sky130_fd_sc_hd__buf_1 _3448_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][0] ),
    .X(_0978_));
 sky130_fd_sc_hd__nor2_2 _3449_ (.A(_0977_),
    .B(_0978_),
    .Y(_0979_));
 sky130_fd_sc_hd__buf_1 _3450_ (.A(_0979_),
    .X(_0980_));
 sky130_fd_sc_hd__buf_1 _3451_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][3] ),
    .X(_0981_));
 sky130_fd_sc_hd__buf_1 _3452_ (.A(_0981_),
    .X(_0982_));
 sky130_fd_sc_hd__buf_1 _3453_ (.A(_0982_),
    .X(_0983_));
 sky130_fd_sc_hd__buf_1 _3454_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][2] ),
    .X(_0984_));
 sky130_fd_sc_hd__buf_1 _3455_ (.A(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__nor2_2 _3456_ (.A(_0983_),
    .B(_0985_),
    .Y(_0986_));
 sky130_fd_sc_hd__nand2_2 _3457_ (.A(_0980_),
    .B(_0986_),
    .Y(_0987_));
 sky130_fd_sc_hd__nor2_2 _3458_ (.A(_0976_),
    .B(_0987_),
    .Y(_0988_));
 sky130_fd_sc_hd__buf_1 _3459_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][8] ),
    .X(_0989_));
 sky130_fd_sc_hd__or2_2 _3460_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][7] ),
    .B(\tree_instances[6].u_tree.pipeline_current_node[0][6] ),
    .X(_0990_));
 sky130_fd_sc_hd__nor2_2 _3461_ (.A(_0989_),
    .B(_0990_),
    .Y(_0991_));
 sky130_fd_sc_hd__a31o_2 _3462_ (.A1(_0971_),
    .A2(_0988_),
    .A3(_0991_),
    .B1(\tree_instances[6].u_tree.tree_state[1] ),
    .X(_0080_));
 sky130_fd_sc_hd__and4_2 _3463_ (.A(\tree_instances[3].u_tree.ready_for_next ),
    .B(\tree_instances[2].u_tree.ready_for_next ),
    .C(\tree_instances[5].u_tree.ready_for_next ),
    .D(\tree_instances[4].u_tree.ready_for_next ),
    .X(_0992_));
 sky130_fd_sc_hd__nand3_2 _3464_ (.A(\tree_instances[1].u_tree.ready_for_next ),
    .B(\tree_instances[0].u_tree.ready_for_next ),
    .C(_0992_),
    .Y(_0993_));
 sky130_fd_sc_hd__and4_2 _3465_ (.A(\tree_instances[11].u_tree.ready_for_next ),
    .B(\tree_instances[10].u_tree.ready_for_next ),
    .C(\tree_instances[13].u_tree.ready_for_next ),
    .D(\tree_instances[12].u_tree.ready_for_next ),
    .X(_0994_));
 sky130_fd_sc_hd__and4_2 _3466_ (.A(\tree_instances[7].u_tree.ready_for_next ),
    .B(\tree_instances[6].u_tree.ready_for_next ),
    .C(\tree_instances[9].u_tree.ready_for_next ),
    .D(\tree_instances[8].u_tree.ready_for_next ),
    .X(_0995_));
 sky130_fd_sc_hd__nand2_2 _3467_ (.A(_0994_),
    .B(_0995_),
    .Y(_0996_));
 sky130_fd_sc_hd__and4_2 _3468_ (.A(\tree_instances[15].u_tree.ready_for_next ),
    .B(\tree_instances[14].u_tree.ready_for_next ),
    .C(\tree_instances[17].u_tree.ready_for_next ),
    .D(\tree_instances[16].u_tree.ready_for_next ),
    .X(_0997_));
 sky130_fd_sc_hd__nand4_2 _3469_ (.A(\tree_instances[19].u_tree.ready_for_next ),
    .B(\tree_instances[18].u_tree.ready_for_next ),
    .C(\tree_instances[20].u_tree.ready_for_next ),
    .D(_0997_),
    .Y(_0998_));
 sky130_fd_sc_hd__nor3_2 _3470_ (.A(_0993_),
    .B(_0996_),
    .C(_0998_),
    .Y(ready_for_next));
 sky130_fd_sc_hd__or2_2 _3471_ (.A(_0731_),
    .B(\tree_instances[8].u_tree.pipeline_valid[0] ),
    .X(_0999_));
 sky130_fd_sc_hd__buf_1 _3472_ (.A(\tree_instances[8].u_tree.tree_state[3] ),
    .X(_1000_));
 sky130_fd_sc_hd__a21o_2 _3473_ (.A1(\tree_instances[8].u_tree.tree_state[0] ),
    .A2(_0999_),
    .B1(_1000_),
    .X(_0083_));
 sky130_fd_sc_hd__buf_1 _3474_ (.A(\tree_instances[7].u_tree.tree_state[2] ),
    .X(_1001_));
 sky130_fd_sc_hd__buf_1 _3475_ (.A(\tree_instances[7].u_tree.pipeline_current_node[0][4] ),
    .X(_1002_));
 sky130_fd_sc_hd__buf_1 _3476_ (.A(\tree_instances[7].u_tree.pipeline_current_node[0][5] ),
    .X(_1003_));
 sky130_fd_sc_hd__or2_2 _3477_ (.A(_1002_),
    .B(_1003_),
    .X(_1004_));
 sky130_fd_sc_hd__buf_1 _3478_ (.A(_1004_),
    .X(_1005_));
 sky130_fd_sc_hd__buf_1 _3479_ (.A(\tree_instances[7].u_tree.pipeline_current_node[0][6] ),
    .X(_1006_));
 sky130_fd_sc_hd__or2_2 _3480_ (.A(_1006_),
    .B(\tree_instances[7].u_tree.pipeline_current_node[0][7] ),
    .X(_1007_));
 sky130_fd_sc_hd__nor2_2 _3481_ (.A(_1005_),
    .B(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__buf_1 _3482_ (.A(\tree_instances[7].u_tree.pipeline_current_node[0][3] ),
    .X(_1009_));
 sky130_fd_sc_hd__or2_2 _3483_ (.A(_1009_),
    .B(\tree_instances[7].u_tree.pipeline_current_node[0][2] ),
    .X(_1010_));
 sky130_fd_sc_hd__buf_1 _3484_ (.A(_1010_),
    .X(_1011_));
 sky130_fd_sc_hd__buf_1 _3485_ (.A(_1011_),
    .X(_1012_));
 sky130_fd_sc_hd__buf_1 _3486_ (.A(\tree_instances[7].u_tree.pipeline_current_node[0][1] ),
    .X(_1013_));
 sky130_fd_sc_hd__buf_1 _3487_ (.A(\tree_instances[7].u_tree.pipeline_current_node[0][0] ),
    .X(_1014_));
 sky130_fd_sc_hd__or2_2 _3488_ (.A(_1013_),
    .B(_1014_),
    .X(_1015_));
 sky130_fd_sc_hd__buf_1 _3489_ (.A(_1015_),
    .X(_1016_));
 sky130_fd_sc_hd__nor2_2 _3490_ (.A(_1012_),
    .B(_1016_),
    .Y(_1017_));
 sky130_fd_sc_hd__a31o_2 _3491_ (.A1(_1001_),
    .A2(_1008_),
    .A3(_1017_),
    .B1(\tree_instances[7].u_tree.tree_state[1] ),
    .X(_0082_));
 sky130_fd_sc_hd__inv_2 _3492_ (.A(\state[1] ),
    .Y(_1018_));
 sky130_fd_sc_hd__or2_2 _3493_ (.A(\state[0] ),
    .B(_1018_),
    .X(_1019_));
 sky130_fd_sc_hd__buf_1 _3494_ (.A(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__inv_2 _3495_ (.A(_1020_),
    .Y(_1021_));
 sky130_fd_sc_hd__buf_1 _3496_ (.A(_1021_),
    .X(_0000_));
 sky130_fd_sc_hd__or2_2 _3497_ (.A(_0732_),
    .B(\tree_instances[16].u_tree.pipeline_valid[0] ),
    .X(_1022_));
 sky130_fd_sc_hd__buf_1 _3498_ (.A(\tree_instances[16].u_tree.tree_state[3] ),
    .X(_1023_));
 sky130_fd_sc_hd__a21o_2 _3499_ (.A1(\tree_instances[16].u_tree.tree_state[0] ),
    .A2(_1022_),
    .B1(_1023_),
    .X(_0059_));
 sky130_fd_sc_hd__or2_2 _3500_ (.A(_0733_),
    .B(\tree_instances[9].u_tree.pipeline_valid[0] ),
    .X(_1024_));
 sky130_fd_sc_hd__buf_1 _3501_ (.A(\tree_instances[9].u_tree.tree_state[3] ),
    .X(_1025_));
 sky130_fd_sc_hd__a21o_2 _3502_ (.A1(\tree_instances[9].u_tree.tree_state[0] ),
    .A2(_1024_),
    .B1(_1025_),
    .X(_0085_));
 sky130_fd_sc_hd__buf_1 _3503_ (.A(\tree_instances[12].u_tree.tree_state[2] ),
    .X(_1026_));
 sky130_fd_sc_hd__buf_1 _3504_ (.A(_0833_),
    .X(_1027_));
 sky130_fd_sc_hd__buf_1 _3505_ (.A(_1027_),
    .X(_1028_));
 sky130_fd_sc_hd__buf_1 _3506_ (.A(_0843_),
    .X(_1029_));
 sky130_fd_sc_hd__nor2_2 _3507_ (.A(_1028_),
    .B(_1029_),
    .Y(_1030_));
 sky130_fd_sc_hd__buf_1 _3508_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][7] ),
    .X(_1031_));
 sky130_fd_sc_hd__buf_1 _3509_ (.A(_0846_),
    .X(_1032_));
 sky130_fd_sc_hd__nor2_2 _3510_ (.A(_1031_),
    .B(_1032_),
    .Y(_1033_));
 sky130_fd_sc_hd__a31o_2 _3511_ (.A1(_1026_),
    .A2(_1030_),
    .A3(_1033_),
    .B1(\tree_instances[12].u_tree.tree_state[1] ),
    .X(_0052_));
 sky130_fd_sc_hd__buf_1 _3512_ (.A(\tree_instances[8].u_tree.tree_state[2] ),
    .X(_1034_));
 sky130_fd_sc_hd__buf_1 _3513_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][7] ),
    .X(_1035_));
 sky130_fd_sc_hd__buf_1 _3514_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][6] ),
    .X(_1036_));
 sky130_fd_sc_hd__buf_1 _3515_ (.A(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__nor2_2 _3516_ (.A(_1035_),
    .B(_1037_),
    .Y(_1038_));
 sky130_fd_sc_hd__buf_1 _3517_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][0] ),
    .X(_1039_));
 sky130_fd_sc_hd__or2_2 _3518_ (.A(_1039_),
    .B(\tree_instances[8].u_tree.pipeline_current_node[0][3] ),
    .X(_1040_));
 sky130_fd_sc_hd__buf_1 _3519_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][1] ),
    .X(_1041_));
 sky130_fd_sc_hd__buf_1 _3520_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][2] ),
    .X(_1042_));
 sky130_fd_sc_hd__or2_2 _3521_ (.A(_1041_),
    .B(_1042_),
    .X(_1043_));
 sky130_fd_sc_hd__buf_1 _3522_ (.A(_1043_),
    .X(_1044_));
 sky130_fd_sc_hd__nor2_2 _3523_ (.A(_1040_),
    .B(_1044_),
    .Y(_1045_));
 sky130_fd_sc_hd__buf_1 _3524_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][4] ),
    .X(_1046_));
 sky130_fd_sc_hd__buf_1 _3525_ (.A(_1046_),
    .X(_1047_));
 sky130_fd_sc_hd__buf_1 _3526_ (.A(_1047_),
    .X(_1048_));
 sky130_fd_sc_hd__buf_1 _3527_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][5] ),
    .X(_1049_));
 sky130_fd_sc_hd__nor2_2 _3528_ (.A(_1048_),
    .B(_1049_),
    .Y(_1050_));
 sky130_fd_sc_hd__a41o_2 _3529_ (.A1(_1034_),
    .A2(_1038_),
    .A3(_1045_),
    .A4(_1050_),
    .B1(\tree_instances[8].u_tree.tree_state[1] ),
    .X(_0084_));
 sky130_fd_sc_hd__buf_1 _3530_ (.A(\tree_instances[15].u_tree.tree_state[2] ),
    .X(_1051_));
 sky130_fd_sc_hd__buf_1 _3531_ (.A(\tree_instances[15].u_tree.pipeline_current_node[0][7] ),
    .X(_1052_));
 sky130_fd_sc_hd__buf_1 _3532_ (.A(_1052_),
    .X(_1053_));
 sky130_fd_sc_hd__buf_1 _3533_ (.A(\tree_instances[15].u_tree.pipeline_current_node[0][6] ),
    .X(_1054_));
 sky130_fd_sc_hd__or2_2 _3534_ (.A(_1054_),
    .B(\tree_instances[15].u_tree.pipeline_current_node[0][5] ),
    .X(_1055_));
 sky130_fd_sc_hd__buf_1 _3535_ (.A(_1055_),
    .X(_1056_));
 sky130_fd_sc_hd__buf_1 _3536_ (.A(_1056_),
    .X(_1057_));
 sky130_fd_sc_hd__nor2_2 _3537_ (.A(_1053_),
    .B(_1057_),
    .Y(_1058_));
 sky130_fd_sc_hd__buf_1 _3538_ (.A(\tree_instances[15].u_tree.pipeline_current_node[0][0] ),
    .X(_1059_));
 sky130_fd_sc_hd__buf_1 _3539_ (.A(_1059_),
    .X(_1060_));
 sky130_fd_sc_hd__buf_1 _3540_ (.A(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__buf_1 _3541_ (.A(\tree_instances[15].u_tree.pipeline_current_node[0][3] ),
    .X(_1062_));
 sky130_fd_sc_hd__or2_2 _3542_ (.A(_1062_),
    .B(\tree_instances[15].u_tree.pipeline_current_node[0][4] ),
    .X(_1063_));
 sky130_fd_sc_hd__or2_2 _3543_ (.A(_1061_),
    .B(_1063_),
    .X(_1064_));
 sky130_fd_sc_hd__or2_2 _3544_ (.A(\tree_instances[15].u_tree.pipeline_current_node[0][1] ),
    .B(\tree_instances[15].u_tree.pipeline_current_node[0][2] ),
    .X(_1065_));
 sky130_fd_sc_hd__buf_1 _3545_ (.A(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__nor2_2 _3546_ (.A(_1064_),
    .B(_1066_),
    .Y(_1067_));
 sky130_fd_sc_hd__a31o_2 _3547_ (.A1(_1051_),
    .A2(_1058_),
    .A3(_1067_),
    .B1(\tree_instances[15].u_tree.tree_state[1] ),
    .X(_0058_));
 sky130_fd_sc_hd__buf_1 _3548_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][0] ),
    .X(_1068_));
 sky130_fd_sc_hd__buf_1 _3549_ (.A(_1068_),
    .X(_1069_));
 sky130_fd_sc_hd__buf_1 _3550_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][3] ),
    .X(_1070_));
 sky130_fd_sc_hd__or2_2 _3551_ (.A(_1069_),
    .B(_1070_),
    .X(_1071_));
 sky130_fd_sc_hd__buf_1 _3552_ (.A(_1071_),
    .X(_1072_));
 sky130_fd_sc_hd__or2_2 _3553_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][1] ),
    .B(\tree_instances[14].u_tree.pipeline_current_node[0][2] ),
    .X(_1073_));
 sky130_fd_sc_hd__buf_1 _3554_ (.A(_1073_),
    .X(_1074_));
 sky130_fd_sc_hd__or2_2 _3555_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][6] ),
    .B(\tree_instances[14].u_tree.pipeline_current_node[0][7] ),
    .X(_1075_));
 sky130_fd_sc_hd__buf_1 _3556_ (.A(_1075_),
    .X(_1076_));
 sky130_fd_sc_hd__or2_2 _3557_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][4] ),
    .B(\tree_instances[14].u_tree.pipeline_current_node[0][5] ),
    .X(_1077_));
 sky130_fd_sc_hd__buf_1 _3558_ (.A(_1077_),
    .X(_1078_));
 sky130_fd_sc_hd__buf_1 _3559_ (.A(_1078_),
    .X(_1079_));
 sky130_fd_sc_hd__buf_1 _3560_ (.A(\tree_instances[14].u_tree.tree_state[2] ),
    .X(_1080_));
 sky130_fd_sc_hd__o41a_2 _3561_ (.A1(_1072_),
    .A2(_1074_),
    .A3(_1076_),
    .A4(_1079_),
    .B1(_1080_),
    .X(_0013_));
 sky130_fd_sc_hd__nor2_2 _3562_ (.A(_1072_),
    .B(_1074_),
    .Y(_1081_));
 sky130_fd_sc_hd__buf_1 _3563_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][6] ),
    .X(_1082_));
 sky130_fd_sc_hd__buf_1 _3564_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][7] ),
    .X(_1083_));
 sky130_fd_sc_hd__nor2_2 _3565_ (.A(_1082_),
    .B(_1083_),
    .Y(_1084_));
 sky130_fd_sc_hd__buf_1 _3566_ (.A(_1084_),
    .X(_1085_));
 sky130_fd_sc_hd__buf_1 _3567_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][4] ),
    .X(_1086_));
 sky130_fd_sc_hd__buf_1 _3568_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][5] ),
    .X(_1087_));
 sky130_fd_sc_hd__nor2_2 _3569_ (.A(_1086_),
    .B(_1087_),
    .Y(_1088_));
 sky130_fd_sc_hd__buf_1 _3570_ (.A(_1088_),
    .X(_1089_));
 sky130_fd_sc_hd__buf_1 _3571_ (.A(_1089_),
    .X(_1090_));
 sky130_fd_sc_hd__a41o_2 _3572_ (.A1(_1080_),
    .A2(_1081_),
    .A3(_1085_),
    .A4(_1090_),
    .B1(\tree_instances[14].u_tree.tree_state[1] ),
    .X(_0056_));
 sky130_fd_sc_hd__buf_1 _3573_ (.A(\tree_instances[9].u_tree.tree_state[2] ),
    .X(_1091_));
 sky130_fd_sc_hd__buf_1 _3574_ (.A(_1091_),
    .X(_1092_));
 sky130_fd_sc_hd__buf_1 _3575_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][6] ),
    .X(_1093_));
 sky130_fd_sc_hd__buf_1 _3576_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][7] ),
    .X(_1094_));
 sky130_fd_sc_hd__nor2_2 _3577_ (.A(_1093_),
    .B(_1094_),
    .Y(_1095_));
 sky130_fd_sc_hd__buf_1 _3578_ (.A(_1095_),
    .X(_1096_));
 sky130_fd_sc_hd__buf_1 _3579_ (.A(_1096_),
    .X(_1097_));
 sky130_fd_sc_hd__nor2_2 _3580_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][0] ),
    .B(\tree_instances[9].u_tree.pipeline_current_node[0][1] ),
    .Y(_1098_));
 sky130_fd_sc_hd__nor2_2 _3581_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][2] ),
    .B(\tree_instances[9].u_tree.pipeline_current_node[0][3] ),
    .Y(_1099_));
 sky130_fd_sc_hd__nand2_2 _3582_ (.A(_1098_),
    .B(_1099_),
    .Y(_1100_));
 sky130_fd_sc_hd__or2_2 _3583_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][5] ),
    .B(\tree_instances[9].u_tree.pipeline_current_node[0][4] ),
    .X(_1101_));
 sky130_fd_sc_hd__buf_1 _3584_ (.A(_1101_),
    .X(_1102_));
 sky130_fd_sc_hd__buf_1 _3585_ (.A(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__nor2_2 _3586_ (.A(_1100_),
    .B(_1103_),
    .Y(_1104_));
 sky130_fd_sc_hd__a31o_2 _3587_ (.A1(_1092_),
    .A2(_1097_),
    .A3(_1104_),
    .B1(\tree_instances[9].u_tree.tree_state[1] ),
    .X(_0086_));
 sky130_fd_sc_hd__inv_2 _3588_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][7] ),
    .Y(_1105_));
 sky130_fd_sc_hd__nor2_2 _3589_ (.A(_1049_),
    .B(_1036_),
    .Y(_1106_));
 sky130_fd_sc_hd__buf_1 _3590_ (.A(_1106_),
    .X(_1107_));
 sky130_fd_sc_hd__nand2_2 _3591_ (.A(_1105_),
    .B(_1107_),
    .Y(_1108_));
 sky130_fd_sc_hd__inv_2 _3592_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][4] ),
    .Y(_1109_));
 sky130_fd_sc_hd__buf_1 _3593_ (.A(_1109_),
    .X(_1110_));
 sky130_fd_sc_hd__nand2_2 _3594_ (.A(_1110_),
    .B(_1045_),
    .Y(_1111_));
 sky130_fd_sc_hd__o21a_2 _3595_ (.A1(_1108_),
    .A2(_1111_),
    .B1(\tree_instances[8].u_tree.tree_state[2] ),
    .X(_0041_));
 sky130_fd_sc_hd__buf_1 _3596_ (.A(_0730_),
    .X(_1112_));
 sky130_fd_sc_hd__or2_2 _3597_ (.A(_1112_),
    .B(\tree_instances[13].u_tree.pipeline_valid[0] ),
    .X(_1113_));
 sky130_fd_sc_hd__buf_1 _3598_ (.A(\tree_instances[13].u_tree.tree_state[3] ),
    .X(_1114_));
 sky130_fd_sc_hd__a21o_2 _3599_ (.A1(\tree_instances[13].u_tree.tree_state[0] ),
    .A2(_1113_),
    .B1(_1114_),
    .X(_0053_));
 sky130_fd_sc_hd__a21boi_2 _3600_ (.A1(_1058_),
    .A2(_1067_),
    .B1_N(_1051_),
    .Y(_0015_));
 sky130_fd_sc_hd__buf_1 _3601_ (.A(\tree_instances[0].u_tree.tree_state[2] ),
    .X(_1115_));
 sky130_fd_sc_hd__buf_1 _3602_ (.A(\tree_instances[0].u_tree.pipeline_current_node[0][7] ),
    .X(_1116_));
 sky130_fd_sc_hd__buf_1 _3603_ (.A(\tree_instances[0].u_tree.pipeline_current_node[0][5] ),
    .X(_1117_));
 sky130_fd_sc_hd__or2_2 _3604_ (.A(\tree_instances[0].u_tree.pipeline_current_node[0][6] ),
    .B(_1117_),
    .X(_1118_));
 sky130_fd_sc_hd__buf_1 _3605_ (.A(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__nor2_2 _3606_ (.A(_1116_),
    .B(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__buf_1 _3607_ (.A(_1120_),
    .X(_1121_));
 sky130_fd_sc_hd__buf_1 _3608_ (.A(\tree_instances[0].u_tree.pipeline_current_node[0][1] ),
    .X(_1122_));
 sky130_fd_sc_hd__buf_1 _3609_ (.A(_1122_),
    .X(_1123_));
 sky130_fd_sc_hd__buf_1 _3610_ (.A(_1123_),
    .X(_1124_));
 sky130_fd_sc_hd__buf_1 _3611_ (.A(\tree_instances[0].u_tree.pipeline_current_node[0][0] ),
    .X(_1125_));
 sky130_fd_sc_hd__buf_1 _3612_ (.A(\tree_instances[0].u_tree.pipeline_current_node[0][2] ),
    .X(_1126_));
 sky130_fd_sc_hd__buf_1 _3613_ (.A(_1126_),
    .X(_1127_));
 sky130_fd_sc_hd__nor2_2 _3614_ (.A(_1125_),
    .B(_1127_),
    .Y(_1128_));
 sky130_fd_sc_hd__buf_1 _3615_ (.A(\tree_instances[0].u_tree.pipeline_current_node[0][4] ),
    .X(_1129_));
 sky130_fd_sc_hd__buf_1 _3616_ (.A(\tree_instances[0].u_tree.pipeline_current_node[0][3] ),
    .X(_1130_));
 sky130_fd_sc_hd__buf_1 _3617_ (.A(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__nor2_2 _3618_ (.A(_1129_),
    .B(_1131_),
    .Y(_1132_));
 sky130_fd_sc_hd__nand2_2 _3619_ (.A(_1128_),
    .B(_1132_),
    .Y(_1133_));
 sky130_fd_sc_hd__nor2_2 _3620_ (.A(_1124_),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__a31o_2 _3621_ (.A1(_1115_),
    .A2(_1121_),
    .A3(_1134_),
    .B1(\tree_instances[0].u_tree.tree_state[1] ),
    .X(_0046_));
 sky130_fd_sc_hd__a21boi_2 _3622_ (.A1(_1121_),
    .A2(_1134_),
    .B1_N(_1115_),
    .Y(_0003_));
 sky130_fd_sc_hd__or2_2 _3623_ (.A(_0731_),
    .B(\tree_instances[10].u_tree.pipeline_valid[0] ),
    .X(_1135_));
 sky130_fd_sc_hd__buf_1 _3624_ (.A(\tree_instances[10].u_tree.tree_state[3] ),
    .X(_1136_));
 sky130_fd_sc_hd__a21o_2 _3625_ (.A1(\tree_instances[10].u_tree.tree_state[0] ),
    .A2(_1135_),
    .B1(_1136_),
    .X(_0047_));
 sky130_fd_sc_hd__buf_1 _3626_ (.A(\tree_instances[15].u_tree.tree_state[3] ),
    .X(_1137_));
 sky130_fd_sc_hd__o21a_2 _3627_ (.A1(_0732_),
    .A2(\tree_instances[15].u_tree.pipeline_valid[0] ),
    .B1(\tree_instances[15].u_tree.tree_state[0] ),
    .X(_1138_));
 sky130_fd_sc_hd__or2_2 _3628_ (.A(_1137_),
    .B(_1138_),
    .X(_1139_));
 sky130_fd_sc_hd__buf_1 _3629_ (.A(_1139_),
    .X(_0057_));
 sky130_fd_sc_hd__buf_1 _3630_ (.A(\tree_instances[11].u_tree.tree_state[2] ),
    .X(_1140_));
 sky130_fd_sc_hd__buf_1 _3631_ (.A(\tree_instances[11].u_tree.pipeline_current_node[0][4] ),
    .X(_1141_));
 sky130_fd_sc_hd__or2_2 _3632_ (.A(_1141_),
    .B(\tree_instances[11].u_tree.pipeline_current_node[0][5] ),
    .X(_1142_));
 sky130_fd_sc_hd__buf_1 _3633_ (.A(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__buf_1 _3634_ (.A(\tree_instances[11].u_tree.pipeline_current_node[0][0] ),
    .X(_1144_));
 sky130_fd_sc_hd__buf_1 _3635_ (.A(\tree_instances[11].u_tree.pipeline_current_node[0][3] ),
    .X(_1145_));
 sky130_fd_sc_hd__or2_2 _3636_ (.A(_1144_),
    .B(_1145_),
    .X(_1146_));
 sky130_fd_sc_hd__buf_1 _3637_ (.A(_1146_),
    .X(_1147_));
 sky130_fd_sc_hd__nor2_2 _3638_ (.A(_1143_),
    .B(_1147_),
    .Y(_1148_));
 sky130_fd_sc_hd__buf_1 _3639_ (.A(\tree_instances[11].u_tree.pipeline_current_node[0][6] ),
    .X(_1149_));
 sky130_fd_sc_hd__nor2_2 _3640_ (.A(_1149_),
    .B(\tree_instances[11].u_tree.pipeline_current_node[0][7] ),
    .Y(_1150_));
 sky130_fd_sc_hd__buf_1 _3641_ (.A(_1150_),
    .X(_1151_));
 sky130_fd_sc_hd__buf_1 _3642_ (.A(_1151_),
    .X(_1152_));
 sky130_fd_sc_hd__buf_1 _3643_ (.A(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__buf_1 _3644_ (.A(\tree_instances[11].u_tree.pipeline_current_node[0][1] ),
    .X(_1154_));
 sky130_fd_sc_hd__buf_1 _3645_ (.A(\tree_instances[11].u_tree.pipeline_current_node[0][2] ),
    .X(_1155_));
 sky130_fd_sc_hd__nor2_2 _3646_ (.A(_1154_),
    .B(_1155_),
    .Y(_1156_));
 sky130_fd_sc_hd__a41o_2 _3647_ (.A1(_1140_),
    .A2(_1148_),
    .A3(_1153_),
    .A4(_1156_),
    .B1(\tree_instances[11].u_tree.tree_state[1] ),
    .X(_0050_));
 sky130_fd_sc_hd__buf_1 _3648_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][7] ),
    .X(_1157_));
 sky130_fd_sc_hd__or2_2 _3649_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][6] ),
    .B(_1157_),
    .X(_1158_));
 sky130_fd_sc_hd__buf_1 _3650_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][2] ),
    .X(_1159_));
 sky130_fd_sc_hd__or2_2 _3651_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][3] ),
    .B(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__buf_1 _3652_ (.A(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__buf_1 _3653_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][1] ),
    .X(_1162_));
 sky130_fd_sc_hd__or2_2 _3654_ (.A(_1162_),
    .B(\tree_instances[10].u_tree.pipeline_current_node[0][0] ),
    .X(_1163_));
 sky130_fd_sc_hd__buf_1 _3655_ (.A(_1163_),
    .X(_1164_));
 sky130_fd_sc_hd__buf_1 _3656_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][4] ),
    .X(_1165_));
 sky130_fd_sc_hd__or2_2 _3657_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][5] ),
    .B(_1165_),
    .X(_1166_));
 sky130_fd_sc_hd__buf_1 _3658_ (.A(_1166_),
    .X(_1167_));
 sky130_fd_sc_hd__buf_1 _3659_ (.A(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__or4_2 _3660_ (.A(_1158_),
    .B(_1161_),
    .C(_1164_),
    .D(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__nand2_2 _3661_ (.A(\tree_instances[10].u_tree.tree_state[2] ),
    .B(_1169_),
    .Y(_1170_));
 sky130_fd_sc_hd__inv_2 _3662_ (.A(_1170_),
    .Y(_0005_));
 sky130_fd_sc_hd__buf_1 _3663_ (.A(\tree_instances[10].u_tree.tree_state[2] ),
    .X(_1171_));
 sky130_fd_sc_hd__buf_1 _3664_ (.A(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__inv_2 _3665_ (.A(_1169_),
    .Y(_0379_));
 sky130_fd_sc_hd__a21o_2 _3666_ (.A1(_1172_),
    .A2(_0379_),
    .B1(\tree_instances[10].u_tree.tree_state[1] ),
    .X(_0048_));
 sky130_fd_sc_hd__buf_1 _3667_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][4] ),
    .X(_1173_));
 sky130_fd_sc_hd__buf_1 _3668_ (.A(_1173_),
    .X(_1174_));
 sky130_fd_sc_hd__buf_1 _3669_ (.A(_1174_),
    .X(_1175_));
 sky130_fd_sc_hd__buf_1 _3670_ (.A(_1175_),
    .X(_1176_));
 sky130_fd_sc_hd__inv_2 _3671_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][7] ),
    .Y(_1177_));
 sky130_fd_sc_hd__buf_1 _3672_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][5] ),
    .X(_1178_));
 sky130_fd_sc_hd__buf_1 _3673_ (.A(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__nor2_2 _3674_ (.A(_1179_),
    .B(\tree_instances[20].u_tree.pipeline_current_node[0][6] ),
    .Y(_1180_));
 sky130_fd_sc_hd__nand2_2 _3675_ (.A(_1177_),
    .B(_1180_),
    .Y(_1181_));
 sky130_fd_sc_hd__nor2_2 _3676_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][1] ),
    .B(\tree_instances[20].u_tree.pipeline_current_node[0][0] ),
    .Y(_1182_));
 sky130_fd_sc_hd__nor2_2 _3677_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][3] ),
    .B(_0766_),
    .Y(_1183_));
 sky130_fd_sc_hd__nand2_2 _3678_ (.A(_1182_),
    .B(_1183_),
    .Y(_1184_));
 sky130_fd_sc_hd__o31a_2 _3679_ (.A1(_1176_),
    .A2(_1181_),
    .A3(_1184_),
    .B1(_0756_),
    .X(_0027_));
 sky130_fd_sc_hd__or2_2 _3680_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][5] ),
    .B(_0852_),
    .X(_1185_));
 sky130_fd_sc_hd__buf_1 _3681_ (.A(_1185_),
    .X(_1186_));
 sky130_fd_sc_hd__buf_1 _3682_ (.A(_0855_),
    .X(_1187_));
 sky130_fd_sc_hd__buf_1 _3683_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][0] ),
    .X(_1188_));
 sky130_fd_sc_hd__buf_1 _3684_ (.A(_1188_),
    .X(_1189_));
 sky130_fd_sc_hd__nor2_2 _3685_ (.A(_1187_),
    .B(_1189_),
    .Y(_1190_));
 sky130_fd_sc_hd__buf_1 _3686_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][3] ),
    .X(_1191_));
 sky130_fd_sc_hd__buf_1 _3687_ (.A(_0858_),
    .X(_1192_));
 sky130_fd_sc_hd__nor2_2 _3688_ (.A(_1191_),
    .B(_1192_),
    .Y(_1193_));
 sky130_fd_sc_hd__nand2_2 _3689_ (.A(_1190_),
    .B(_1193_),
    .Y(_1194_));
 sky130_fd_sc_hd__buf_1 _3690_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][7] ),
    .X(_1195_));
 sky130_fd_sc_hd__or2_2 _3691_ (.A(_1195_),
    .B(_0862_),
    .X(_1196_));
 sky130_fd_sc_hd__o31a_2 _3692_ (.A1(_1186_),
    .A2(_1194_),
    .A3(_1196_),
    .B1(_0850_),
    .X(_0031_));
 sky130_fd_sc_hd__a21boi_2 _3693_ (.A1(_0809_),
    .A2(_0828_),
    .B1_N(_0802_),
    .Y(_0029_));
 sky130_fd_sc_hd__buf_1 _3694_ (.A(\tree_instances[20].u_tree.tree_state[3] ),
    .X(_1197_));
 sky130_fd_sc_hd__o21ai_2 _3695_ (.A1(_0731_),
    .A2(\tree_instances[20].u_tree.pipeline_valid[0] ),
    .B1(\tree_instances[20].u_tree.tree_state[0] ),
    .Y(_1198_));
 sky130_fd_sc_hd__or2b_2 _3696_ (.A(_1197_),
    .B_N(_1198_),
    .X(_1199_));
 sky130_fd_sc_hd__buf_1 _3697_ (.A(_1199_),
    .X(_0069_));
 sky130_fd_sc_hd__buf_1 _3698_ (.A(_1143_),
    .X(_1200_));
 sky130_fd_sc_hd__buf_1 _3699_ (.A(_1149_),
    .X(_1201_));
 sky130_fd_sc_hd__buf_1 _3700_ (.A(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__buf_1 _3701_ (.A(\tree_instances[11].u_tree.pipeline_current_node[0][7] ),
    .X(_1203_));
 sky130_fd_sc_hd__or2_2 _3702_ (.A(_1202_),
    .B(_1203_),
    .X(_1204_));
 sky130_fd_sc_hd__or2_2 _3703_ (.A(\tree_instances[11].u_tree.pipeline_current_node[0][1] ),
    .B(\tree_instances[11].u_tree.pipeline_current_node[0][2] ),
    .X(_1205_));
 sky130_fd_sc_hd__o41a_2 _3704_ (.A1(_1200_),
    .A2(_1147_),
    .A3(_1204_),
    .A4(_1205_),
    .B1(_1140_),
    .X(_0007_));
 sky130_fd_sc_hd__or2_2 _3705_ (.A(_1093_),
    .B(\tree_instances[9].u_tree.pipeline_current_node[0][7] ),
    .X(_1206_));
 sky130_fd_sc_hd__o31a_2 _3706_ (.A1(_1206_),
    .A2(_1100_),
    .A3(_1103_),
    .B1(_1092_),
    .X(_0043_));
 sky130_fd_sc_hd__buf_1 _3707_ (.A(_1005_),
    .X(_1207_));
 sky130_fd_sc_hd__buf_1 _3708_ (.A(_1007_),
    .X(_1208_));
 sky130_fd_sc_hd__buf_1 _3709_ (.A(\tree_instances[7].u_tree.pipeline_current_node[0][2] ),
    .X(_1209_));
 sky130_fd_sc_hd__nor2_2 _3710_ (.A(_1009_),
    .B(_1209_),
    .Y(_1210_));
 sky130_fd_sc_hd__buf_1 _3711_ (.A(_1210_),
    .X(_1211_));
 sky130_fd_sc_hd__buf_1 _3712_ (.A(_1013_),
    .X(_1212_));
 sky130_fd_sc_hd__nor2_2 _3713_ (.A(_1212_),
    .B(_1014_),
    .Y(_1213_));
 sky130_fd_sc_hd__nand2_2 _3714_ (.A(_1211_),
    .B(_1213_),
    .Y(_1214_));
 sky130_fd_sc_hd__o31a_2 _3715_ (.A1(_1207_),
    .A2(_1208_),
    .A3(_1214_),
    .B1(_1001_),
    .X(_0039_));
 sky130_fd_sc_hd__or2_2 _3716_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][7] ),
    .B(_0914_),
    .X(_1215_));
 sky130_fd_sc_hd__buf_1 _3717_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][1] ),
    .X(_1216_));
 sky130_fd_sc_hd__buf_1 _3718_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][0] ),
    .X(_1217_));
 sky130_fd_sc_hd__nor2_2 _3719_ (.A(_1216_),
    .B(_1217_),
    .Y(_1218_));
 sky130_fd_sc_hd__buf_1 _3720_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][2] ),
    .X(_1219_));
 sky130_fd_sc_hd__nor2_2 _3721_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][3] ),
    .B(_1219_),
    .Y(_1220_));
 sky130_fd_sc_hd__nand2_2 _3722_ (.A(_1218_),
    .B(_1220_),
    .Y(_1221_));
 sky130_fd_sc_hd__buf_1 _3723_ (.A(_0926_),
    .X(_1222_));
 sky130_fd_sc_hd__or2_2 _3724_ (.A(_0925_),
    .B(_1222_),
    .X(_1223_));
 sky130_fd_sc_hd__buf_1 _3725_ (.A(_1223_),
    .X(_1224_));
 sky130_fd_sc_hd__buf_1 _3726_ (.A(_1224_),
    .X(_1225_));
 sky130_fd_sc_hd__o31a_2 _3727_ (.A1(_1215_),
    .A2(_1221_),
    .A3(_1225_),
    .B1(\tree_instances[16].u_tree.tree_state[2] ),
    .X(_0017_));
 sky130_fd_sc_hd__or2_2 _3728_ (.A(_0731_),
    .B(\tree_instances[1].u_tree.pipeline_valid[0] ),
    .X(_1226_));
 sky130_fd_sc_hd__buf_1 _3729_ (.A(\tree_instances[1].u_tree.tree_state[3] ),
    .X(_1227_));
 sky130_fd_sc_hd__a21o_2 _3730_ (.A1(\tree_instances[1].u_tree.tree_state[0] ),
    .A2(_1226_),
    .B1(_1227_),
    .X(_0067_));
 sky130_fd_sc_hd__buf_1 _3731_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][7] ),
    .X(_1228_));
 sky130_fd_sc_hd__buf_1 _3732_ (.A(_0897_),
    .X(_1229_));
 sky130_fd_sc_hd__or2_2 _3733_ (.A(_1229_),
    .B(_0898_),
    .X(_1230_));
 sky130_fd_sc_hd__buf_1 _3734_ (.A(_1230_),
    .X(_1231_));
 sky130_fd_sc_hd__nor2_2 _3735_ (.A(_1228_),
    .B(_1231_),
    .Y(_1232_));
 sky130_fd_sc_hd__a31o_2 _3736_ (.A1(_0901_),
    .A2(_0894_),
    .A3(_1232_),
    .B1(\tree_instances[19].u_tree.tree_state[1] ),
    .X(_0066_));
 sky130_fd_sc_hd__buf_1 _3737_ (.A(_0989_),
    .X(_1233_));
 sky130_fd_sc_hd__buf_1 _3738_ (.A(_0990_),
    .X(_1234_));
 sky130_fd_sc_hd__or2_2 _3739_ (.A(_0976_),
    .B(_0987_),
    .X(_1235_));
 sky130_fd_sc_hd__o31a_2 _3740_ (.A1(_1233_),
    .A2(_1234_),
    .A3(_1235_),
    .B1(_0971_),
    .X(_0037_));
 sky130_fd_sc_hd__or2_2 _3741_ (.A(_0792_),
    .B(_0793_),
    .X(_1236_));
 sky130_fd_sc_hd__buf_1 _3742_ (.A(_1236_),
    .X(_1237_));
 sky130_fd_sc_hd__buf_1 _3743_ (.A(_0791_),
    .X(_1238_));
 sky130_fd_sc_hd__nand2_2 _3744_ (.A(_1238_),
    .B(_0777_),
    .Y(_1239_));
 sky130_fd_sc_hd__o31a_2 _3745_ (.A1(_0789_),
    .A2(_1237_),
    .A3(_1239_),
    .B1(_0776_),
    .X(_0019_));
 sky130_fd_sc_hd__buf_1 _3746_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][0] ),
    .X(_1240_));
 sky130_fd_sc_hd__nor2_2 _3747_ (.A(_1240_),
    .B(\tree_instances[5].u_tree.pipeline_current_node[0][1] ),
    .Y(_1241_));
 sky130_fd_sc_hd__buf_1 _3748_ (.A(_1241_),
    .X(_1242_));
 sky130_fd_sc_hd__nor2_2 _3749_ (.A(_0937_),
    .B(_0939_),
    .Y(_1243_));
 sky130_fd_sc_hd__buf_1 _3750_ (.A(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__nand2_2 _3751_ (.A(_1242_),
    .B(_1244_),
    .Y(_1245_));
 sky130_fd_sc_hd__or2_2 _3752_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][7] ),
    .B(_0945_),
    .X(_1246_));
 sky130_fd_sc_hd__inv_2 _3753_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][6] ),
    .Y(_1247_));
 sky130_fd_sc_hd__buf_1 _3754_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][4] ),
    .X(_1248_));
 sky130_fd_sc_hd__nor2_2 _3755_ (.A(_1248_),
    .B(\tree_instances[5].u_tree.pipeline_current_node[0][5] ),
    .Y(_1249_));
 sky130_fd_sc_hd__nand2_2 _3756_ (.A(_1247_),
    .B(_1249_),
    .Y(_1250_));
 sky130_fd_sc_hd__o31a_2 _3757_ (.A1(_1245_),
    .A2(_1246_),
    .A3(_1250_),
    .B1(\tree_instances[5].u_tree.tree_state[2] ),
    .X(_0035_));
 sky130_fd_sc_hd__or2_2 _3758_ (.A(_0732_),
    .B(\tree_instances[19].u_tree.pipeline_valid[0] ),
    .X(_1251_));
 sky130_fd_sc_hd__buf_1 _3759_ (.A(\tree_instances[19].u_tree.tree_state[3] ),
    .X(_1252_));
 sky130_fd_sc_hd__a21o_2 _3760_ (.A1(\tree_instances[19].u_tree.tree_state[0] ),
    .A2(_1251_),
    .B1(_1252_),
    .X(_0065_));
 sky130_fd_sc_hd__buf_1 _3761_ (.A(_0746_),
    .X(_1253_));
 sky130_fd_sc_hd__nor2_2 _3762_ (.A(_1253_),
    .B(_0742_),
    .Y(_1254_));
 sky130_fd_sc_hd__buf_1 _3763_ (.A(_0745_),
    .X(_1255_));
 sky130_fd_sc_hd__buf_1 _3764_ (.A(_1255_),
    .X(_1256_));
 sky130_fd_sc_hd__buf_1 _3765_ (.A(_1256_),
    .X(_1257_));
 sky130_fd_sc_hd__nor2_2 _3766_ (.A(_1257_),
    .B(_0744_),
    .Y(_1258_));
 sky130_fd_sc_hd__a31o_2 _3767_ (.A1(_0751_),
    .A2(_1254_),
    .A3(_1258_),
    .B1(\tree_instances[18].u_tree.tree_state[1] ),
    .X(_0064_));
 sky130_fd_sc_hd__and2b_2 _3768_ (.A_N(\tree_instances[7].u_tree.prediction_valid ),
    .B(_0970_),
    .X(_1259_));
 sky130_fd_sc_hd__buf_1 _3769_ (.A(_1259_),
    .X(_0105_));
 sky130_fd_sc_hd__buf_1 _3770_ (.A(_1144_),
    .X(_1260_));
 sky130_fd_sc_hd__buf_1 _3771_ (.A(_1260_),
    .X(_1261_));
 sky130_fd_sc_hd__buf_1 _3772_ (.A(\tree_instances[11].u_tree.pipeline_current_node[0][2] ),
    .X(_1262_));
 sky130_fd_sc_hd__buf_1 _3773_ (.A(_1145_),
    .X(_1263_));
 sky130_fd_sc_hd__buf_1 _3774_ (.A(_1263_),
    .X(_1264_));
 sky130_fd_sc_hd__buf_1 _3775_ (.A(_1264_),
    .X(_1265_));
 sky130_fd_sc_hd__buf_1 _3776_ (.A(_1154_),
    .X(_1266_));
 sky130_fd_sc_hd__buf_1 _3777_ (.A(_1141_),
    .X(_1267_));
 sky130_fd_sc_hd__buf_1 _3778_ (.A(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__buf_1 _3779_ (.A(\tree_instances[11].u_tree.pipeline_current_node[0][5] ),
    .X(_1269_));
 sky130_fd_sc_hd__buf_1 _3780_ (.A(_1265_),
    .X(_1270_));
 sky130_fd_sc_hd__buf_1 _3781_ (.A(_1270_),
    .X(_1271_));
 sky130_fd_sc_hd__buf_1 _3782_ (.A(_1262_),
    .X(_1272_));
 sky130_fd_sc_hd__buf_1 _3783_ (.A(_1272_),
    .X(_1273_));
 sky130_fd_sc_hd__buf_1 _3784_ (.A(_1273_),
    .X(_1274_));
 sky130_fd_sc_hd__buf_1 _3785_ (.A(_1261_),
    .X(_1275_));
 sky130_fd_sc_hd__buf_1 _3786_ (.A(_1266_),
    .X(_1276_));
 sky130_fd_sc_hd__buf_1 _3787_ (.A(_1268_),
    .X(_1277_));
 sky130_fd_sc_hd__buf_1 _3788_ (.A(_1271_),
    .X(_1278_));
 sky130_fd_sc_hd__buf_1 _3789_ (.A(_1269_),
    .X(_1279_));
 sky130_fd_sc_hd__buf_1 _3790_ (.A(_1279_),
    .X(_1280_));
 sky130_fd_sc_hd__buf_1 _3791_ (.A(_1280_),
    .X(_1281_));
 sky130_fd_sc_hd__buf_1 _3792_ (.A(_1277_),
    .X(_1282_));
 sky130_fd_sc_hd__buf_1 _3793_ (.A(_1201_),
    .X(_1283_));
 sky130_fd_sc_hd__buf_1 _3794_ (.A(_1282_),
    .X(_1284_));
 sky130_fd_sc_hd__buf_1 _3795_ (.A(_1203_),
    .X(_1285_));
 sky130_fd_sc_hd__buf_1 _3796_ (.A(_1283_),
    .X(_1286_));
 sky130_fd_sc_hd__and2b_2 _3797_ (.A_N(\tree_instances[8].u_tree.prediction_valid ),
    .B(_1000_),
    .X(_1287_));
 sky130_fd_sc_hd__buf_1 _3798_ (.A(_1287_),
    .X(_0106_));
 sky130_fd_sc_hd__buf_1 _3799_ (.A(\tree_instances[7].u_tree.pipeline_current_node[0][7] ),
    .X(_1288_));
 sky130_fd_sc_hd__buf_1 _3800_ (.A(_1014_),
    .X(_1289_));
 sky130_fd_sc_hd__buf_1 _3801_ (.A(_1289_),
    .X(_1290_));
 sky130_fd_sc_hd__buf_1 _3802_ (.A(_1212_),
    .X(_1291_));
 sky130_fd_sc_hd__buf_1 _3803_ (.A(_1209_),
    .X(_1292_));
 sky130_fd_sc_hd__buf_1 _3804_ (.A(_1003_),
    .X(_1293_));
 sky130_fd_sc_hd__buf_1 _3805_ (.A(_1002_),
    .X(_1294_));
 sky130_fd_sc_hd__buf_1 _3806_ (.A(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__buf_1 _3807_ (.A(_1295_),
    .X(_1296_));
 sky130_fd_sc_hd__buf_1 _3808_ (.A(_1296_),
    .X(_1297_));
 sky130_fd_sc_hd__buf_1 _3809_ (.A(_1288_),
    .X(_1298_));
 sky130_fd_sc_hd__buf_1 _3810_ (.A(_1293_),
    .X(_1299_));
 sky130_fd_sc_hd__buf_1 _3811_ (.A(_1299_),
    .X(_1300_));
 sky130_fd_sc_hd__buf_1 _3812_ (.A(_1298_),
    .X(_1301_));
 sky130_fd_sc_hd__buf_1 _3813_ (.A(_1301_),
    .X(_1302_));
 sky130_fd_sc_hd__buf_1 _3814_ (.A(_1291_),
    .X(_1303_));
 sky130_fd_sc_hd__buf_1 _3815_ (.A(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__buf_1 _3816_ (.A(_1297_),
    .X(_1305_));
 sky130_fd_sc_hd__buf_1 _3817_ (.A(_1009_),
    .X(_1306_));
 sky130_fd_sc_hd__buf_1 _3818_ (.A(_1306_),
    .X(_1307_));
 sky130_fd_sc_hd__buf_1 _3819_ (.A(_1307_),
    .X(_1308_));
 sky130_fd_sc_hd__buf_1 _3820_ (.A(_1308_),
    .X(_1309_));
 sky130_fd_sc_hd__buf_1 _3821_ (.A(_1292_),
    .X(_1310_));
 sky130_fd_sc_hd__buf_1 _3822_ (.A(_1006_),
    .X(_1311_));
 sky130_fd_sc_hd__buf_1 _3823_ (.A(_1311_),
    .X(_1312_));
 sky130_fd_sc_hd__buf_1 _3824_ (.A(_1312_),
    .X(_1313_));
 sky130_fd_sc_hd__and2b_2 _3825_ (.A_N(\tree_instances[9].u_tree.prediction_valid ),
    .B(_1025_),
    .X(_1314_));
 sky130_fd_sc_hd__buf_1 _3826_ (.A(_1314_),
    .X(_0107_));
 sky130_fd_sc_hd__and2b_2 _3827_ (.A_N(\tree_instances[10].u_tree.prediction_valid ),
    .B(_1136_),
    .X(_1315_));
 sky130_fd_sc_hd__buf_1 _3828_ (.A(_1315_),
    .X(_0088_));
 sky130_fd_sc_hd__nor2_2 _3829_ (.A(_0951_),
    .B(\tree_instances[11].u_tree.prediction_valid ),
    .Y(_0089_));
 sky130_fd_sc_hd__and2b_2 _3830_ (.A_N(\tree_instances[12].u_tree.prediction_valid ),
    .B(_0829_),
    .X(_1316_));
 sky130_fd_sc_hd__buf_1 _3831_ (.A(_1316_),
    .X(_0090_));
 sky130_fd_sc_hd__buf_1 _3832_ (.A(_1195_),
    .X(_1317_));
 sky130_fd_sc_hd__buf_1 _3833_ (.A(_1191_),
    .X(_1318_));
 sky130_fd_sc_hd__inv_2 _3834_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][4] ),
    .Y(_1319_));
 sky130_fd_sc_hd__buf_1 _3835_ (.A(_1189_),
    .X(_1320_));
 sky130_fd_sc_hd__buf_1 _3836_ (.A(_1318_),
    .X(_1321_));
 sky130_fd_sc_hd__inv_2 _3837_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][1] ),
    .Y(_1322_));
 sky130_fd_sc_hd__buf_1 _3838_ (.A(_0858_),
    .X(_1323_));
 sky130_fd_sc_hd__buf_1 _3839_ (.A(_0852_),
    .X(_1324_));
 sky130_fd_sc_hd__buf_1 _3840_ (.A(_1320_),
    .X(_1325_));
 sky130_fd_sc_hd__buf_1 _3841_ (.A(_0862_),
    .X(_1326_));
 sky130_fd_sc_hd__buf_1 _3842_ (.A(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__inv_2 _3843_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][3] ),
    .Y(_1328_));
 sky130_fd_sc_hd__buf_1 _3844_ (.A(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__buf_1 _3845_ (.A(_1187_),
    .X(_1330_));
 sky130_fd_sc_hd__buf_1 _3846_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][5] ),
    .X(_1331_));
 sky130_fd_sc_hd__buf_1 _3847_ (.A(_1192_),
    .X(_1332_));
 sky130_fd_sc_hd__buf_1 _3848_ (.A(_1324_),
    .X(_1333_));
 sky130_fd_sc_hd__buf_1 _3849_ (.A(_1333_),
    .X(_1334_));
 sky130_fd_sc_hd__inv_2 _3850_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][6] ),
    .Y(_1335_));
 sky130_fd_sc_hd__and2b_2 _3851_ (.A_N(_1188_),
    .B(\tree_instances[3].u_tree.pipeline_current_node[0][3] ),
    .X(_1336_));
 sky130_fd_sc_hd__nor2_2 _3852_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][5] ),
    .B(\tree_instances[3].u_tree.pipeline_current_node[0][6] ),
    .Y(_1337_));
 sky130_fd_sc_hd__buf_1 _3853_ (.A(_1332_),
    .X(_1338_));
 sky130_fd_sc_hd__and2_2 _3854_ (.A(_1187_),
    .B(_1323_),
    .X(_1339_));
 sky130_fd_sc_hd__nand2_2 _3855_ (.A(_1339_),
    .B(_1336_),
    .Y(_1340_));
 sky130_fd_sc_hd__buf_1 _3856_ (.A(_1334_),
    .X(_1341_));
 sky130_fd_sc_hd__buf_1 _3857_ (.A(_1331_),
    .X(_1342_));
 sky130_fd_sc_hd__buf_1 _3858_ (.A(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__buf_1 _3859_ (.A(_1341_),
    .X(_1344_));
 sky130_fd_sc_hd__buf_1 _3860_ (.A(_1317_),
    .X(_1345_));
 sky130_fd_sc_hd__buf_1 _3861_ (.A(_1345_),
    .X(_1346_));
 sky130_fd_sc_hd__buf_1 _3862_ (.A(_1321_),
    .X(_1347_));
 sky130_fd_sc_hd__nor2_2 _3863_ (.A(_1324_),
    .B(_1340_),
    .Y(_1348_));
 sky130_fd_sc_hd__and3_2 _3864_ (.A(_1195_),
    .B(_1337_),
    .C(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__buf_1 _3865_ (.A(_1349_),
    .X(_0489_));
 sky130_fd_sc_hd__buf_1 _3866_ (.A(_1338_),
    .X(_1350_));
 sky130_fd_sc_hd__buf_1 _3867_ (.A(_1330_),
    .X(_1351_));
 sky130_fd_sc_hd__buf_1 _3868_ (.A(_1343_),
    .X(_1352_));
 sky130_fd_sc_hd__inv_2 _3869_ (.A(_1217_),
    .Y(_1353_));
 sky130_fd_sc_hd__buf_1 _3870_ (.A(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__inv_2 _3871_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][3] ),
    .Y(_1355_));
 sky130_fd_sc_hd__nor2_2 _3872_ (.A(_1355_),
    .B(_0926_),
    .Y(_1356_));
 sky130_fd_sc_hd__nor2b_2 _3873_ (.A(_1219_),
    .B_N(_1216_),
    .Y(_1357_));
 sky130_fd_sc_hd__nand2_2 _3874_ (.A(_1356_),
    .B(_1357_),
    .Y(_1358_));
 sky130_fd_sc_hd__nor2_2 _3875_ (.A(_1354_),
    .B(_1358_),
    .Y(_1359_));
 sky130_fd_sc_hd__buf_1 _3876_ (.A(_0925_),
    .X(_1360_));
 sky130_fd_sc_hd__buf_1 _3877_ (.A(_1360_),
    .X(_1361_));
 sky130_fd_sc_hd__nand2_2 _3878_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][7] ),
    .B(\tree_instances[16].u_tree.pipeline_current_node[0][6] ),
    .Y(_1362_));
 sky130_fd_sc_hd__nor2_2 _3879_ (.A(_1361_),
    .B(_1362_),
    .Y(_1363_));
 sky130_fd_sc_hd__a32o_2 _3880_ (.A1(_0918_),
    .A2(_0924_),
    .A3(_0930_),
    .B1(_1359_),
    .B2(_1363_),
    .X(_0001_));
 sky130_fd_sc_hd__buf_1 _3881_ (.A(_1222_),
    .X(_1364_));
 sky130_fd_sc_hd__buf_1 _3882_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][0] ),
    .X(_1365_));
 sky130_fd_sc_hd__buf_1 _3883_ (.A(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__buf_1 _3884_ (.A(_1216_),
    .X(_1367_));
 sky130_fd_sc_hd__inv_2 _3885_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][7] ),
    .Y(_1368_));
 sky130_fd_sc_hd__buf_1 _3886_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][3] ),
    .X(_1369_));
 sky130_fd_sc_hd__buf_1 _3887_ (.A(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__buf_1 _3888_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][2] ),
    .X(_1371_));
 sky130_fd_sc_hd__buf_1 _3889_ (.A(_1364_),
    .X(_1372_));
 sky130_fd_sc_hd__buf_1 _3890_ (.A(_1372_),
    .X(_1373_));
 sky130_fd_sc_hd__buf_1 _3891_ (.A(_1360_),
    .X(_1374_));
 sky130_fd_sc_hd__buf_1 _3892_ (.A(_1219_),
    .X(_1375_));
 sky130_fd_sc_hd__buf_1 _3893_ (.A(_0913_),
    .X(_1376_));
 sky130_fd_sc_hd__buf_1 _3894_ (.A(_1370_),
    .X(_1377_));
 sky130_fd_sc_hd__buf_1 _3895_ (.A(_1371_),
    .X(_1378_));
 sky130_fd_sc_hd__buf_1 _3896_ (.A(_1367_),
    .X(_1379_));
 sky130_fd_sc_hd__buf_1 _3897_ (.A(_1373_),
    .X(_1380_));
 sky130_fd_sc_hd__buf_1 _3898_ (.A(_1374_),
    .X(_1381_));
 sky130_fd_sc_hd__buf_1 _3899_ (.A(_1378_),
    .X(_1382_));
 sky130_fd_sc_hd__buf_1 _3900_ (.A(_1381_),
    .X(_1383_));
 sky130_fd_sc_hd__buf_1 _3901_ (.A(_1377_),
    .X(_1384_));
 sky130_fd_sc_hd__buf_1 _3902_ (.A(_0913_),
    .X(_1385_));
 sky130_fd_sc_hd__buf_1 _3903_ (.A(_1366_),
    .X(_1386_));
 sky130_fd_sc_hd__buf_1 _3904_ (.A(_0915_),
    .X(_1387_));
 sky130_fd_sc_hd__buf_1 _3905_ (.A(_1387_),
    .X(_1388_));
 sky130_fd_sc_hd__and2b_2 _3906_ (.A_N(\tree_instances[13].u_tree.prediction_valid ),
    .B(_1114_),
    .X(_1389_));
 sky130_fd_sc_hd__buf_1 _3907_ (.A(_1389_),
    .X(_0091_));
 sky130_fd_sc_hd__and2b_2 _3908_ (.A_N(\tree_instances[14].u_tree.prediction_valid ),
    .B(_0735_),
    .X(_1390_));
 sky130_fd_sc_hd__buf_1 _3909_ (.A(_1390_),
    .X(_0092_));
 sky130_fd_sc_hd__and2b_2 _3910_ (.A_N(\tree_instances[15].u_tree.prediction_valid ),
    .B(_1137_),
    .X(_1391_));
 sky130_fd_sc_hd__buf_1 _3911_ (.A(_1391_),
    .X(_0093_));
 sky130_fd_sc_hd__buf_1 _3912_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][7] ),
    .X(_1392_));
 sky130_fd_sc_hd__inv_2 _3913_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][6] ),
    .Y(_1393_));
 sky130_fd_sc_hd__buf_1 _3914_ (.A(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__inv_2 _3915_ (.A(_1173_),
    .Y(_1395_));
 sky130_fd_sc_hd__buf_1 _3916_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][1] ),
    .X(_1396_));
 sky130_fd_sc_hd__buf_1 _3917_ (.A(_1396_),
    .X(_1397_));
 sky130_fd_sc_hd__buf_1 _3918_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][2] ),
    .X(_1398_));
 sky130_fd_sc_hd__inv_2 _3919_ (.A(_1398_),
    .Y(_1399_));
 sky130_fd_sc_hd__buf_1 _3920_ (.A(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__buf_1 _3921_ (.A(_1183_),
    .X(_1401_));
 sky130_fd_sc_hd__inv_2 _3922_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][3] ),
    .Y(_1402_));
 sky130_fd_sc_hd__buf_1 _3923_ (.A(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__buf_1 _3924_ (.A(_1397_),
    .X(_1404_));
 sky130_fd_sc_hd__buf_1 _3925_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][0] ),
    .X(_1405_));
 sky130_fd_sc_hd__buf_1 _3926_ (.A(_1405_),
    .X(_1406_));
 sky130_fd_sc_hd__buf_1 _3927_ (.A(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__buf_1 _3928_ (.A(_0758_),
    .X(_1408_));
 sky130_fd_sc_hd__inv_2 _3929_ (.A(\tree_instances[20].u_tree.pipeline_current_node[0][0] ),
    .Y(_1409_));
 sky130_fd_sc_hd__buf_1 _3930_ (.A(_1409_),
    .X(_1410_));
 sky130_fd_sc_hd__buf_1 _3931_ (.A(_1404_),
    .X(_1411_));
 sky130_fd_sc_hd__nor2_2 _3932_ (.A(_1177_),
    .B(_1394_),
    .Y(_1412_));
 sky130_fd_sc_hd__buf_1 _3933_ (.A(_0764_),
    .X(_1413_));
 sky130_fd_sc_hd__buf_1 _3934_ (.A(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__buf_1 _3935_ (.A(_1414_),
    .X(_1415_));
 sky130_fd_sc_hd__and2_2 _3936_ (.A(_1397_),
    .B(_1409_),
    .X(_1416_));
 sky130_fd_sc_hd__buf_1 _3937_ (.A(_1392_),
    .X(_1417_));
 sky130_fd_sc_hd__buf_1 _3938_ (.A(_1417_),
    .X(_1418_));
 sky130_fd_sc_hd__buf_1 _3939_ (.A(_1408_),
    .X(_1419_));
 sky130_fd_sc_hd__buf_1 _3940_ (.A(_1176_),
    .X(_1420_));
 sky130_fd_sc_hd__buf_1 _3941_ (.A(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__buf_1 _3942_ (.A(_1411_),
    .X(_1422_));
 sky130_fd_sc_hd__buf_1 _3943_ (.A(_1179_),
    .X(_1423_));
 sky130_fd_sc_hd__buf_1 _3944_ (.A(_1423_),
    .X(_1424_));
 sky130_fd_sc_hd__buf_1 _3945_ (.A(_1417_),
    .X(_1425_));
 sky130_fd_sc_hd__buf_1 _3946_ (.A(_1416_),
    .X(_1426_));
 sky130_fd_sc_hd__buf_1 _3947_ (.A(_0758_),
    .X(_1427_));
 sky130_fd_sc_hd__buf_1 _3948_ (.A(_1427_),
    .X(_1428_));
 sky130_fd_sc_hd__buf_1 _3949_ (.A(_1412_),
    .X(_1429_));
 sky130_fd_sc_hd__and3_2 _3950_ (.A(_1401_),
    .B(_0771_),
    .C(_1426_),
    .X(_1430_));
 sky130_fd_sc_hd__buf_1 _3951_ (.A(_0767_),
    .X(_1431_));
 sky130_fd_sc_hd__buf_1 _3952_ (.A(_1415_),
    .X(_1432_));
 sky130_fd_sc_hd__buf_1 _3953_ (.A(_1419_),
    .X(_1433_));
 sky130_fd_sc_hd__buf_1 _3954_ (.A(\tree_instances[15].u_tree.pipeline_current_node[0][2] ),
    .X(_1434_));
 sky130_fd_sc_hd__buf_1 _3955_ (.A(\tree_instances[15].u_tree.pipeline_current_node[0][4] ),
    .X(_1435_));
 sky130_fd_sc_hd__buf_1 _3956_ (.A(\tree_instances[15].u_tree.pipeline_current_node[0][1] ),
    .X(_1436_));
 sky130_fd_sc_hd__buf_1 _3957_ (.A(\tree_instances[15].u_tree.pipeline_current_node[0][5] ),
    .X(_1437_));
 sky130_fd_sc_hd__buf_1 _3958_ (.A(_1434_),
    .X(_1438_));
 sky130_fd_sc_hd__buf_1 _3959_ (.A(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__buf_1 _3960_ (.A(_1435_),
    .X(_1440_));
 sky130_fd_sc_hd__buf_1 _3961_ (.A(_1061_),
    .X(_1441_));
 sky130_fd_sc_hd__buf_1 _3962_ (.A(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__buf_1 _3963_ (.A(_1052_),
    .X(_1443_));
 sky130_fd_sc_hd__buf_1 _3964_ (.A(_1443_),
    .X(_1444_));
 sky130_fd_sc_hd__buf_1 _3965_ (.A(_1440_),
    .X(_1445_));
 sky130_fd_sc_hd__buf_1 _3966_ (.A(_1437_),
    .X(_1446_));
 sky130_fd_sc_hd__buf_1 _3967_ (.A(_1062_),
    .X(_1447_));
 sky130_fd_sc_hd__buf_1 _3968_ (.A(_1054_),
    .X(_1448_));
 sky130_fd_sc_hd__buf_1 _3969_ (.A(_1445_),
    .X(_1449_));
 sky130_fd_sc_hd__buf_1 _3970_ (.A(_1447_),
    .X(_1450_));
 sky130_fd_sc_hd__buf_1 _3971_ (.A(_1448_),
    .X(_1451_));
 sky130_fd_sc_hd__buf_1 _3972_ (.A(_1446_),
    .X(_1452_));
 sky130_fd_sc_hd__buf_1 _3973_ (.A(_1452_),
    .X(_1453_));
 sky130_fd_sc_hd__buf_1 _3974_ (.A(_1439_),
    .X(_1454_));
 sky130_fd_sc_hd__buf_1 _3975_ (.A(_1436_),
    .X(_1455_));
 sky130_fd_sc_hd__buf_1 _3976_ (.A(_1449_),
    .X(_1456_));
 sky130_fd_sc_hd__buf_1 _3977_ (.A(_1450_),
    .X(_1457_));
 sky130_fd_sc_hd__and2b_2 _3978_ (.A_N(\tree_instances[16].u_tree.prediction_valid ),
    .B(_1023_),
    .X(_1458_));
 sky130_fd_sc_hd__buf_1 _3979_ (.A(_1458_),
    .X(_0094_));
 sky130_fd_sc_hd__inv_2 _3980_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][7] ),
    .Y(_1459_));
 sky130_fd_sc_hd__buf_1 _3981_ (.A(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__inv_2 _3982_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][6] ),
    .Y(_1461_));
 sky130_fd_sc_hd__nor2_2 _3983_ (.A(_1460_),
    .B(_1461_),
    .Y(_1462_));
 sky130_fd_sc_hd__buf_1 _3984_ (.A(_1462_),
    .X(_1463_));
 sky130_fd_sc_hd__buf_1 _3985_ (.A(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__inv_2 _3986_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][5] ),
    .Y(_1465_));
 sky130_fd_sc_hd__buf_1 _3987_ (.A(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__buf_1 _3988_ (.A(_1466_),
    .X(_1467_));
 sky130_fd_sc_hd__buf_1 _3989_ (.A(_1467_),
    .X(_1468_));
 sky130_fd_sc_hd__buf_1 _3990_ (.A(_0868_),
    .X(_1469_));
 sky130_fd_sc_hd__nor2_2 _3991_ (.A(_1469_),
    .B(_0877_),
    .Y(_1470_));
 sky130_fd_sc_hd__inv_2 _3992_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][2] ),
    .Y(_1471_));
 sky130_fd_sc_hd__nand2_2 _3993_ (.A(_0867_),
    .B(_0870_),
    .Y(_1472_));
 sky130_fd_sc_hd__nor2_2 _3994_ (.A(_1471_),
    .B(_1472_),
    .Y(_1473_));
 sky130_fd_sc_hd__nand2_2 _3995_ (.A(_1470_),
    .B(_1473_),
    .Y(_1474_));
 sky130_fd_sc_hd__nor2_2 _3996_ (.A(_1468_),
    .B(_1474_),
    .Y(_1475_));
 sky130_fd_sc_hd__a21o_2 _3997_ (.A1(_1464_),
    .A2(_1475_),
    .B1(_0883_),
    .X(_0002_));
 sky130_fd_sc_hd__buf_1 _3998_ (.A(_0877_),
    .X(_1476_));
 sky130_fd_sc_hd__buf_1 _3999_ (.A(_0879_),
    .X(_1477_));
 sky130_fd_sc_hd__buf_1 _4000_ (.A(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__buf_1 _4001_ (.A(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__buf_1 _4002_ (.A(_1479_),
    .X(_1480_));
 sky130_fd_sc_hd__buf_1 _4003_ (.A(_1471_),
    .X(_1481_));
 sky130_fd_sc_hd__buf_1 _4004_ (.A(_0871_),
    .X(_1482_));
 sky130_fd_sc_hd__buf_1 _4005_ (.A(\tree_instances[1].u_tree.pipeline_current_node[0][6] ),
    .X(_1483_));
 sky130_fd_sc_hd__buf_1 _4006_ (.A(_1469_),
    .X(_1484_));
 sky130_fd_sc_hd__buf_1 _4007_ (.A(_1484_),
    .X(_1485_));
 sky130_fd_sc_hd__buf_1 _4008_ (.A(_1476_),
    .X(_1486_));
 sky130_fd_sc_hd__buf_1 _4009_ (.A(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__buf_1 _4010_ (.A(_0867_),
    .X(_1488_));
 sky130_fd_sc_hd__buf_1 _4011_ (.A(_1483_),
    .X(_1489_));
 sky130_fd_sc_hd__buf_1 _4012_ (.A(_0876_),
    .X(_1490_));
 sky130_fd_sc_hd__buf_1 _4013_ (.A(_0872_),
    .X(_1491_));
 sky130_fd_sc_hd__buf_1 _4014_ (.A(_1488_),
    .X(_1492_));
 sky130_fd_sc_hd__buf_1 _4015_ (.A(_1485_),
    .X(_1493_));
 sky130_fd_sc_hd__buf_1 _4016_ (.A(_1491_),
    .X(_1494_));
 sky130_fd_sc_hd__buf_1 _4017_ (.A(_1487_),
    .X(_1495_));
 sky130_fd_sc_hd__buf_1 _4018_ (.A(_1482_),
    .X(_1496_));
 sky130_fd_sc_hd__buf_1 _4019_ (.A(_1493_),
    .X(_1497_));
 sky130_fd_sc_hd__buf_1 _4020_ (.A(_1490_),
    .X(_1498_));
 sky130_fd_sc_hd__and2b_2 _4021_ (.A_N(\tree_instances[17].u_tree.prediction_valid ),
    .B(_0909_),
    .X(_1499_));
 sky130_fd_sc_hd__buf_1 _4022_ (.A(_1499_),
    .X(_0095_));
 sky130_fd_sc_hd__buf_1 _4023_ (.A(_0885_),
    .X(_1500_));
 sky130_fd_sc_hd__buf_1 _4024_ (.A(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__buf_1 _4025_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][0] ),
    .X(_1502_));
 sky130_fd_sc_hd__buf_1 _4026_ (.A(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__buf_1 _4027_ (.A(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__buf_1 _4028_ (.A(\tree_instances[19].u_tree.pipeline_current_node[0][1] ),
    .X(_1505_));
 sky130_fd_sc_hd__buf_1 _4029_ (.A(_0884_),
    .X(_1506_));
 sky130_fd_sc_hd__buf_1 _4030_ (.A(_0898_),
    .X(_1507_));
 sky130_fd_sc_hd__buf_1 _4031_ (.A(_1507_),
    .X(_1508_));
 sky130_fd_sc_hd__buf_1 _4032_ (.A(_1508_),
    .X(_1509_));
 sky130_fd_sc_hd__buf_1 _4033_ (.A(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__buf_1 _4034_ (.A(_1501_),
    .X(_1511_));
 sky130_fd_sc_hd__buf_1 _4035_ (.A(_1505_),
    .X(_1512_));
 sky130_fd_sc_hd__buf_1 _4036_ (.A(_0891_),
    .X(_1513_));
 sky130_fd_sc_hd__buf_1 _4037_ (.A(_1506_),
    .X(_1514_));
 sky130_fd_sc_hd__buf_1 _4038_ (.A(_1513_),
    .X(_1515_));
 sky130_fd_sc_hd__buf_1 _4039_ (.A(_1515_),
    .X(_1516_));
 sky130_fd_sc_hd__buf_1 _4040_ (.A(_1514_),
    .X(_1517_));
 sky130_fd_sc_hd__buf_1 _4041_ (.A(_1229_),
    .X(_1518_));
 sky130_fd_sc_hd__buf_1 _4042_ (.A(_1517_),
    .X(_1519_));
 sky130_fd_sc_hd__buf_1 _4043_ (.A(_1511_),
    .X(_1520_));
 sky130_fd_sc_hd__buf_1 _4044_ (.A(_1228_),
    .X(_1521_));
 sky130_fd_sc_hd__buf_1 _4045_ (.A(_1521_),
    .X(_1522_));
 sky130_fd_sc_hd__buf_1 _4046_ (.A(_1518_),
    .X(_1523_));
 sky130_fd_sc_hd__buf_1 _4047_ (.A(_1523_),
    .X(_1524_));
 sky130_fd_sc_hd__buf_1 _4048_ (.A(_1524_),
    .X(_1525_));
 sky130_fd_sc_hd__buf_1 _4049_ (.A(_1520_),
    .X(_1526_));
 sky130_fd_sc_hd__buf_1 _4050_ (.A(_1504_),
    .X(_1527_));
 sky130_fd_sc_hd__and2b_2 _4051_ (.A_N(\tree_instances[18].u_tree.prediction_valid ),
    .B(_0753_),
    .X(_1528_));
 sky130_fd_sc_hd__buf_1 _4052_ (.A(_1528_),
    .X(_0096_));
 sky130_fd_sc_hd__buf_1 _4053_ (.A(_1070_),
    .X(_1529_));
 sky130_fd_sc_hd__buf_1 _4054_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][1] ),
    .X(_1530_));
 sky130_fd_sc_hd__buf_1 _4055_ (.A(_1069_),
    .X(_1531_));
 sky130_fd_sc_hd__buf_1 _4056_ (.A(\tree_instances[14].u_tree.pipeline_current_node[0][2] ),
    .X(_1532_));
 sky130_fd_sc_hd__buf_1 _4057_ (.A(_1087_),
    .X(_1533_));
 sky130_fd_sc_hd__buf_1 _4058_ (.A(_1531_),
    .X(_1534_));
 sky130_fd_sc_hd__buf_1 _4059_ (.A(_1086_),
    .X(_1535_));
 sky130_fd_sc_hd__buf_1 _4060_ (.A(_1535_),
    .X(_1536_));
 sky130_fd_sc_hd__buf_1 _4061_ (.A(_1530_),
    .X(_1537_));
 sky130_fd_sc_hd__buf_1 _4062_ (.A(_1532_),
    .X(_1538_));
 sky130_fd_sc_hd__buf_1 _4063_ (.A(_1529_),
    .X(_1539_));
 sky130_fd_sc_hd__buf_1 _4064_ (.A(_1539_),
    .X(_1540_));
 sky130_fd_sc_hd__buf_1 _4065_ (.A(_1533_),
    .X(_1541_));
 sky130_fd_sc_hd__buf_1 _4066_ (.A(_1538_),
    .X(_1542_));
 sky130_fd_sc_hd__buf_1 _4067_ (.A(_1541_),
    .X(_1543_));
 sky130_fd_sc_hd__buf_1 _4068_ (.A(_1540_),
    .X(_1544_));
 sky130_fd_sc_hd__buf_1 _4069_ (.A(_1536_),
    .X(_1545_));
 sky130_fd_sc_hd__buf_1 _4070_ (.A(_1537_),
    .X(_1546_));
 sky130_fd_sc_hd__buf_1 _4071_ (.A(_1545_),
    .X(_1547_));
 sky130_fd_sc_hd__and2b_2 _4072_ (.A_N(\tree_instances[19].u_tree.prediction_valid ),
    .B(_1252_),
    .X(_1548_));
 sky130_fd_sc_hd__buf_1 _4073_ (.A(_1548_),
    .X(_0097_));
 sky130_fd_sc_hd__buf_1 _4074_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][6] ),
    .X(_1549_));
 sky130_fd_sc_hd__buf_1 _4075_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][1] ),
    .X(_1550_));
 sky130_fd_sc_hd__buf_1 _4076_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][0] ),
    .X(_1551_));
 sky130_fd_sc_hd__buf_1 _4077_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][2] ),
    .X(_1552_));
 sky130_fd_sc_hd__buf_1 _4078_ (.A(_1551_),
    .X(_1553_));
 sky130_fd_sc_hd__buf_1 _4079_ (.A(\tree_instances[18].u_tree.pipeline_current_node[0][3] ),
    .X(_1554_));
 sky130_fd_sc_hd__buf_1 _4080_ (.A(_1554_),
    .X(_1555_));
 sky130_fd_sc_hd__buf_1 _4081_ (.A(_1555_),
    .X(_1556_));
 sky130_fd_sc_hd__buf_1 _4082_ (.A(_1556_),
    .X(_1557_));
 sky130_fd_sc_hd__buf_1 _4083_ (.A(_0746_),
    .X(_1558_));
 sky130_fd_sc_hd__buf_1 _4084_ (.A(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__buf_1 _4085_ (.A(_0743_),
    .X(_1560_));
 sky130_fd_sc_hd__buf_1 _4086_ (.A(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__buf_1 _4087_ (.A(_1549_),
    .X(_1562_));
 sky130_fd_sc_hd__buf_1 _4088_ (.A(_1562_),
    .X(_1563_));
 sky130_fd_sc_hd__buf_1 _4089_ (.A(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__buf_1 _4090_ (.A(_1559_),
    .X(_1565_));
 sky130_fd_sc_hd__buf_1 _4091_ (.A(_1557_),
    .X(_1566_));
 sky130_fd_sc_hd__buf_1 _4092_ (.A(_1552_),
    .X(_1567_));
 sky130_fd_sc_hd__buf_1 _4093_ (.A(_1553_),
    .X(_1568_));
 sky130_fd_sc_hd__buf_1 _4094_ (.A(_1256_),
    .X(_1569_));
 sky130_fd_sc_hd__buf_1 _4095_ (.A(_1565_),
    .X(_1570_));
 sky130_fd_sc_hd__buf_1 _4096_ (.A(_1550_),
    .X(_1571_));
 sky130_fd_sc_hd__buf_1 _4097_ (.A(_1567_),
    .X(_1572_));
 sky130_fd_sc_hd__buf_1 _4098_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][6] ),
    .X(_1573_));
 sky130_fd_sc_hd__buf_1 _4099_ (.A(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__inv_2 _4100_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][4] ),
    .Y(_1575_));
 sky130_fd_sc_hd__buf_1 _4101_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][3] ),
    .X(_1576_));
 sky130_fd_sc_hd__buf_1 _4102_ (.A(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__inv_2 _4103_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][0] ),
    .Y(_1578_));
 sky130_fd_sc_hd__buf_1 _4104_ (.A(_1578_),
    .X(_1579_));
 sky130_fd_sc_hd__inv_2 _4105_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][1] ),
    .Y(_1580_));
 sky130_fd_sc_hd__buf_1 _4106_ (.A(_1580_),
    .X(_1581_));
 sky130_fd_sc_hd__buf_1 _4107_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][0] ),
    .X(_1582_));
 sky130_fd_sc_hd__buf_1 _4108_ (.A(_1582_),
    .X(_1583_));
 sky130_fd_sc_hd__buf_1 _4109_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][5] ),
    .X(_1584_));
 sky130_fd_sc_hd__buf_1 _4110_ (.A(_1584_),
    .X(_1585_));
 sky130_fd_sc_hd__buf_1 _4111_ (.A(_1575_),
    .X(_1586_));
 sky130_fd_sc_hd__buf_1 _4112_ (.A(_1165_),
    .X(_1587_));
 sky130_fd_sc_hd__buf_1 _4113_ (.A(_1587_),
    .X(_1588_));
 sky130_fd_sc_hd__buf_1 _4114_ (.A(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__buf_1 _4115_ (.A(_1583_),
    .X(_1590_));
 sky130_fd_sc_hd__buf_1 _4116_ (.A(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__buf_1 _4117_ (.A(_1577_),
    .X(_1592_));
 sky130_fd_sc_hd__buf_1 _4118_ (.A(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__buf_1 _4119_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][2] ),
    .X(_1594_));
 sky130_fd_sc_hd__inv_2 _4120_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][6] ),
    .Y(_1595_));
 sky130_fd_sc_hd__inv_2 _4121_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][7] ),
    .Y(_1596_));
 sky130_fd_sc_hd__buf_1 _4122_ (.A(_1162_),
    .X(_1597_));
 sky130_fd_sc_hd__inv_2 _4123_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][3] ),
    .Y(_1598_));
 sky130_fd_sc_hd__buf_1 _4124_ (.A(_1598_),
    .X(_1599_));
 sky130_fd_sc_hd__buf_1 _4125_ (.A(_1594_),
    .X(_1600_));
 sky130_fd_sc_hd__buf_1 _4126_ (.A(_1574_),
    .X(_1601_));
 sky130_fd_sc_hd__buf_1 _4127_ (.A(_1585_),
    .X(_1602_));
 sky130_fd_sc_hd__buf_1 _4128_ (.A(_1157_),
    .X(_1603_));
 sky130_fd_sc_hd__buf_1 _4129_ (.A(_1603_),
    .X(_1604_));
 sky130_fd_sc_hd__buf_1 _4130_ (.A(_1597_),
    .X(_1605_));
 sky130_fd_sc_hd__buf_1 _4131_ (.A(_1599_),
    .X(_1606_));
 sky130_fd_sc_hd__buf_1 _4132_ (.A(_1605_),
    .X(_1607_));
 sky130_fd_sc_hd__buf_1 _4133_ (.A(_1589_),
    .X(_1608_));
 sky130_fd_sc_hd__buf_1 _4134_ (.A(_1587_),
    .X(_1609_));
 sky130_fd_sc_hd__buf_1 _4135_ (.A(_1601_),
    .X(_1610_));
 sky130_fd_sc_hd__buf_1 _4136_ (.A(_1600_),
    .X(_1611_));
 sky130_fd_sc_hd__buf_1 _4137_ (.A(_1602_),
    .X(_1612_));
 sky130_fd_sc_hd__buf_1 _4138_ (.A(_1611_),
    .X(_1613_));
 sky130_fd_sc_hd__buf_1 _4139_ (.A(_1612_),
    .X(_1614_));
 sky130_fd_sc_hd__buf_1 _4140_ (.A(_1593_),
    .X(_1615_));
 sky130_fd_sc_hd__and2b_2 _4141_ (.A_N(\tree_instances[20].u_tree.prediction_valid ),
    .B(_1197_),
    .X(_1616_));
 sky130_fd_sc_hd__buf_1 _4142_ (.A(_1616_),
    .X(_0099_));
 sky130_fd_sc_hd__and2b_2 _4143_ (.A_N(\tree_instances[0].u_tree.prediction_valid ),
    .B(_0737_),
    .X(_1617_));
 sky130_fd_sc_hd__buf_1 _4144_ (.A(_1617_),
    .X(_0087_));
 sky130_fd_sc_hd__and2b_2 _4145_ (.A_N(\tree_instances[1].u_tree.prediction_valid ),
    .B(_1227_),
    .X(_1618_));
 sky130_fd_sc_hd__buf_1 _4146_ (.A(_1618_),
    .X(_0098_));
 sky130_fd_sc_hd__buf_1 _4147_ (.A(\tree_instances[0].u_tree.pipeline_current_node[0][6] ),
    .X(_1619_));
 sky130_fd_sc_hd__buf_1 _4148_ (.A(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__buf_1 _4149_ (.A(_1117_),
    .X(_1621_));
 sky130_fd_sc_hd__buf_1 _4150_ (.A(_1621_),
    .X(_1622_));
 sky130_fd_sc_hd__buf_1 _4151_ (.A(_1622_),
    .X(_1623_));
 sky130_fd_sc_hd__buf_1 _4152_ (.A(_1131_),
    .X(_1624_));
 sky130_fd_sc_hd__buf_1 _4153_ (.A(_1125_),
    .X(_1625_));
 sky130_fd_sc_hd__buf_1 _4154_ (.A(\tree_instances[0].u_tree.pipeline_current_node[0][4] ),
    .X(_1626_));
 sky130_fd_sc_hd__buf_1 _4155_ (.A(_1625_),
    .X(_1627_));
 sky130_fd_sc_hd__buf_1 _4156_ (.A(_1620_),
    .X(_1628_));
 sky130_fd_sc_hd__buf_1 _4157_ (.A(_1127_),
    .X(_1629_));
 sky130_fd_sc_hd__buf_1 _4158_ (.A(_1626_),
    .X(_1630_));
 sky130_fd_sc_hd__buf_1 _4159_ (.A(_1630_),
    .X(_1631_));
 sky130_fd_sc_hd__buf_1 _4160_ (.A(_1116_),
    .X(_1632_));
 sky130_fd_sc_hd__buf_1 _4161_ (.A(_1624_),
    .X(_1633_));
 sky130_fd_sc_hd__buf_1 _4162_ (.A(_1632_),
    .X(_1634_));
 sky130_fd_sc_hd__buf_1 _4163_ (.A(_1629_),
    .X(_1635_));
 sky130_fd_sc_hd__buf_1 _4164_ (.A(_1628_),
    .X(_1636_));
 sky130_fd_sc_hd__buf_1 _4165_ (.A(_1124_),
    .X(_1637_));
 sky130_fd_sc_hd__buf_1 _4166_ (.A(_1635_),
    .X(_1638_));
 sky130_fd_sc_hd__buf_1 _4167_ (.A(_1631_),
    .X(_1639_));
 sky130_fd_sc_hd__inv_2 _4168_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][5] ),
    .Y(_1640_));
 sky130_fd_sc_hd__buf_1 _4169_ (.A(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__buf_1 _4170_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][4] ),
    .X(_1642_));
 sky130_fd_sc_hd__buf_1 _4171_ (.A(_1642_),
    .X(_1643_));
 sky130_fd_sc_hd__buf_1 _4172_ (.A(_1643_),
    .X(_1644_));
 sky130_fd_sc_hd__buf_1 _4173_ (.A(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__buf_1 _4174_ (.A(_1645_),
    .X(_1646_));
 sky130_fd_sc_hd__buf_1 _4175_ (.A(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__buf_1 _4176_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][3] ),
    .X(_1648_));
 sky130_fd_sc_hd__buf_1 _4177_ (.A(_1648_),
    .X(_1649_));
 sky130_fd_sc_hd__buf_1 _4178_ (.A(_1649_),
    .X(_1650_));
 sky130_fd_sc_hd__buf_1 _4179_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][1] ),
    .X(_1651_));
 sky130_fd_sc_hd__buf_1 _4180_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][0] ),
    .X(_1652_));
 sky130_fd_sc_hd__inv_2 _4181_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][2] ),
    .Y(_1653_));
 sky130_fd_sc_hd__buf_1 _4182_ (.A(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__buf_1 _4183_ (.A(_1650_),
    .X(_1655_));
 sky130_fd_sc_hd__inv_2 _4184_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][0] ),
    .Y(_1656_));
 sky130_fd_sc_hd__buf_1 _4185_ (.A(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__buf_1 _4186_ (.A(_0957_),
    .X(_1658_));
 sky130_fd_sc_hd__buf_1 _4187_ (.A(_1652_),
    .X(_1659_));
 sky130_fd_sc_hd__buf_1 _4188_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][5] ),
    .X(_1660_));
 sky130_fd_sc_hd__buf_1 _4189_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][6] ),
    .X(_1661_));
 sky130_fd_sc_hd__inv_2 _4190_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][6] ),
    .Y(_1662_));
 sky130_fd_sc_hd__buf_1 _4191_ (.A(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__buf_1 _4192_ (.A(_1659_),
    .X(_1664_));
 sky130_fd_sc_hd__nor2b_2 _4193_ (.A(_1651_),
    .B_N(_0956_),
    .Y(_1665_));
 sky130_fd_sc_hd__buf_1 _4194_ (.A(_1664_),
    .X(_1666_));
 sky130_fd_sc_hd__buf_1 _4195_ (.A(_1660_),
    .X(_1667_));
 sky130_fd_sc_hd__buf_1 _4196_ (.A(_1661_),
    .X(_1668_));
 sky130_fd_sc_hd__buf_1 _4197_ (.A(_1668_),
    .X(_1669_));
 sky130_fd_sc_hd__nand2_2 _4198_ (.A(_1657_),
    .B(_1665_),
    .Y(_1670_));
 sky130_fd_sc_hd__buf_1 _4199_ (.A(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__buf_1 _4200_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][7] ),
    .X(_1672_));
 sky130_fd_sc_hd__buf_1 _4201_ (.A(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__buf_1 _4202_ (.A(_1667_),
    .X(_1674_));
 sky130_fd_sc_hd__buf_1 _4203_ (.A(_1674_),
    .X(_1675_));
 sky130_fd_sc_hd__buf_1 _4204_ (.A(_1675_),
    .X(_1676_));
 sky130_fd_sc_hd__buf_1 _4205_ (.A(_1655_),
    .X(_1677_));
 sky130_fd_sc_hd__buf_1 _4206_ (.A(_1658_),
    .X(_1678_));
 sky130_fd_sc_hd__buf_1 _4207_ (.A(_1651_),
    .X(_1679_));
 sky130_fd_sc_hd__nor2_2 _4208_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][5] ),
    .B(_1663_),
    .Y(_1680_));
 sky130_fd_sc_hd__or2_2 _4209_ (.A(_1648_),
    .B(\tree_instances[13].u_tree.pipeline_current_node[0][4] ),
    .X(_1681_));
 sky130_fd_sc_hd__buf_1 _4210_ (.A(_1681_),
    .X(_1682_));
 sky130_fd_sc_hd__buf_1 _4211_ (.A(_1680_),
    .X(_1683_));
 sky130_fd_sc_hd__buf_1 _4212_ (.A(_1677_),
    .X(_1684_));
 sky130_fd_sc_hd__nor2_2 _4213_ (.A(_1682_),
    .B(_1671_),
    .Y(_1685_));
 sky130_fd_sc_hd__buf_1 _4214_ (.A(_1678_),
    .X(_1686_));
 sky130_fd_sc_hd__and2b_2 _4215_ (.A_N(\tree_instances[2].u_tree.prediction_valid ),
    .B(_0755_),
    .X(_1687_));
 sky130_fd_sc_hd__buf_1 _4216_ (.A(_1687_),
    .X(_0100_));
 sky130_fd_sc_hd__and2b_2 _4217_ (.A_N(\tree_instances[3].u_tree.prediction_valid ),
    .B(_0799_),
    .X(_1688_));
 sky130_fd_sc_hd__buf_1 _4218_ (.A(_1688_),
    .X(_0101_));
 sky130_fd_sc_hd__and2b_2 _4219_ (.A_N(\tree_instances[4].u_tree.prediction_valid ),
    .B(_0849_),
    .X(_1689_));
 sky130_fd_sc_hd__buf_1 _4220_ (.A(_1689_),
    .X(_0102_));
 sky130_fd_sc_hd__buf_1 _4221_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][4] ),
    .X(_1690_));
 sky130_fd_sc_hd__inv_2 _4222_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][5] ),
    .Y(_1691_));
 sky130_fd_sc_hd__buf_1 _4223_ (.A(_1691_),
    .X(_1692_));
 sky130_fd_sc_hd__buf_1 _4224_ (.A(_1690_),
    .X(_1693_));
 sky130_fd_sc_hd__buf_1 _4225_ (.A(_1693_),
    .X(_1694_));
 sky130_fd_sc_hd__buf_1 _4226_ (.A(_1694_),
    .X(_1695_));
 sky130_fd_sc_hd__buf_1 _4227_ (.A(_1695_),
    .X(_1696_));
 sky130_fd_sc_hd__buf_1 _4228_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][3] ),
    .X(_1697_));
 sky130_fd_sc_hd__inv_2 _4229_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][3] ),
    .Y(_1698_));
 sky130_fd_sc_hd__buf_1 _4230_ (.A(_0834_),
    .X(_1699_));
 sky130_fd_sc_hd__nor2_2 _4231_ (.A(_1692_),
    .B(_1694_),
    .Y(_1700_));
 sky130_fd_sc_hd__buf_1 _4232_ (.A(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__inv_2 _4233_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][0] ),
    .Y(_1702_));
 sky130_fd_sc_hd__buf_1 _4234_ (.A(_0838_),
    .X(_1703_));
 sky130_fd_sc_hd__buf_1 _4235_ (.A(_0840_),
    .X(_1704_));
 sky130_fd_sc_hd__and2b_2 _4236_ (.A_N(_0839_),
    .B(_0837_),
    .X(_1705_));
 sky130_fd_sc_hd__buf_1 _4237_ (.A(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__buf_1 _4238_ (.A(_1699_),
    .X(_1707_));
 sky130_fd_sc_hd__buf_1 _4239_ (.A(_1707_),
    .X(_1708_));
 sky130_fd_sc_hd__inv_2 _4240_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][7] ),
    .Y(_1709_));
 sky130_fd_sc_hd__buf_1 _4241_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][5] ),
    .X(_1710_));
 sky130_fd_sc_hd__inv_2 _4242_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][4] ),
    .Y(_1711_));
 sky130_fd_sc_hd__inv_2 _4243_ (.A(_0845_),
    .Y(_1712_));
 sky130_fd_sc_hd__buf_1 _4244_ (.A(_1703_),
    .X(_1713_));
 sky130_fd_sc_hd__buf_1 _4245_ (.A(_1697_),
    .X(_1714_));
 sky130_fd_sc_hd__buf_1 _4246_ (.A(_1714_),
    .X(_1715_));
 sky130_fd_sc_hd__buf_1 _4247_ (.A(_1715_),
    .X(_1716_));
 sky130_fd_sc_hd__buf_1 _4248_ (.A(_1031_),
    .X(_1717_));
 sky130_fd_sc_hd__buf_1 _4249_ (.A(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__buf_1 _4250_ (.A(_1710_),
    .X(_1719_));
 sky130_fd_sc_hd__buf_1 _4251_ (.A(_1719_),
    .X(_1720_));
 sky130_fd_sc_hd__buf_1 _4252_ (.A(_1720_),
    .X(_1721_));
 sky130_fd_sc_hd__nor2_2 _4253_ (.A(_1709_),
    .B(_1712_),
    .Y(_1722_));
 sky130_fd_sc_hd__buf_1 _4254_ (.A(_1704_),
    .X(_1723_));
 sky130_fd_sc_hd__buf_1 _4255_ (.A(_1716_),
    .X(_1724_));
 sky130_fd_sc_hd__buf_1 _4256_ (.A(_1032_),
    .X(_1725_));
 sky130_fd_sc_hd__buf_1 _4257_ (.A(_1725_),
    .X(_1726_));
 sky130_fd_sc_hd__buf_1 _4258_ (.A(_1696_),
    .X(_1727_));
 sky130_fd_sc_hd__and2b_2 _4259_ (.A_N(\tree_instances[5].u_tree.prediction_valid ),
    .B(_0903_),
    .X(_1728_));
 sky130_fd_sc_hd__buf_1 _4260_ (.A(_1728_),
    .X(_0103_));
 sky130_fd_sc_hd__buf_1 _4261_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][4] ),
    .X(_1729_));
 sky130_fd_sc_hd__buf_1 _4262_ (.A(_1729_),
    .X(_1730_));
 sky130_fd_sc_hd__buf_1 _4263_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][0] ),
    .X(_1731_));
 sky130_fd_sc_hd__buf_1 _4264_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][1] ),
    .X(_1732_));
 sky130_fd_sc_hd__buf_1 _4265_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][2] ),
    .X(_1733_));
 sky130_fd_sc_hd__buf_1 _4266_ (.A(_1733_),
    .X(_1734_));
 sky130_fd_sc_hd__buf_1 _4267_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][3] ),
    .X(_1735_));
 sky130_fd_sc_hd__buf_1 _4268_ (.A(_1735_),
    .X(_1736_));
 sky130_fd_sc_hd__buf_1 _4269_ (.A(\tree_instances[9].u_tree.pipeline_current_node[0][5] ),
    .X(_1737_));
 sky130_fd_sc_hd__buf_1 _4270_ (.A(_1737_),
    .X(_1738_));
 sky130_fd_sc_hd__buf_1 _4271_ (.A(_1732_),
    .X(_1739_));
 sky130_fd_sc_hd__buf_1 _4272_ (.A(_1738_),
    .X(_1740_));
 sky130_fd_sc_hd__buf_1 _4273_ (.A(_1739_),
    .X(_1741_));
 sky130_fd_sc_hd__buf_1 _4274_ (.A(_1741_),
    .X(_1742_));
 sky130_fd_sc_hd__buf_1 _4275_ (.A(_1731_),
    .X(_1743_));
 sky130_fd_sc_hd__buf_1 _4276_ (.A(_1730_),
    .X(_1744_));
 sky130_fd_sc_hd__buf_1 _4277_ (.A(_1744_),
    .X(_1745_));
 sky130_fd_sc_hd__buf_1 _4278_ (.A(_1736_),
    .X(_1746_));
 sky130_fd_sc_hd__buf_1 _4279_ (.A(_1746_),
    .X(_1747_));
 sky130_fd_sc_hd__buf_1 _4280_ (.A(_1740_),
    .X(_1748_));
 sky130_fd_sc_hd__buf_1 _4281_ (.A(_1748_),
    .X(_1749_));
 sky130_fd_sc_hd__buf_1 _4282_ (.A(_1743_),
    .X(_1750_));
 sky130_fd_sc_hd__buf_1 _4283_ (.A(_1094_),
    .X(_1751_));
 sky130_fd_sc_hd__buf_1 _4284_ (.A(_1751_),
    .X(_1752_));
 sky130_fd_sc_hd__buf_1 _4285_ (.A(_1093_),
    .X(_1753_));
 sky130_fd_sc_hd__buf_1 _4286_ (.A(_1753_),
    .X(_1754_));
 sky130_fd_sc_hd__buf_1 _4287_ (.A(_1754_),
    .X(_1755_));
 sky130_fd_sc_hd__buf_1 _4288_ (.A(_1747_),
    .X(_1756_));
 sky130_fd_sc_hd__buf_1 _4289_ (.A(_1756_),
    .X(_1757_));
 sky130_fd_sc_hd__buf_1 _4290_ (.A(_1745_),
    .X(_1758_));
 sky130_fd_sc_hd__buf_1 _4291_ (.A(_1758_),
    .X(_1759_));
 sky130_fd_sc_hd__buf_1 _4292_ (.A(_1734_),
    .X(_1760_));
 sky130_fd_sc_hd__and2b_2 _4293_ (.A_N(\tree_instances[6].u_tree.prediction_valid ),
    .B(_0932_),
    .X(_1761_));
 sky130_fd_sc_hd__buf_1 _4294_ (.A(_1761_),
    .X(_0104_));
 sky130_fd_sc_hd__buf_1 _4295_ (.A(_1037_),
    .X(_1762_));
 sky130_fd_sc_hd__buf_1 _4296_ (.A(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__buf_1 _4297_ (.A(_1763_),
    .X(_1764_));
 sky130_fd_sc_hd__buf_1 _4298_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][3] ),
    .X(_1765_));
 sky130_fd_sc_hd__nand2b_2 _4299_ (.A_N(\tree_instances[8].u_tree.pipeline_current_node[0][0] ),
    .B(\tree_instances[8].u_tree.pipeline_current_node[0][2] ),
    .Y(_1766_));
 sky130_fd_sc_hd__or2_2 _4300_ (.A(_1041_),
    .B(_1766_),
    .X(_1767_));
 sky130_fd_sc_hd__buf_1 _4301_ (.A(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__buf_1 _4302_ (.A(_1042_),
    .X(_1769_));
 sky130_fd_sc_hd__buf_1 _4303_ (.A(_1765_),
    .X(_1770_));
 sky130_fd_sc_hd__buf_1 _4304_ (.A(_1769_),
    .X(_1771_));
 sky130_fd_sc_hd__inv_2 _4305_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][3] ),
    .Y(_1772_));
 sky130_fd_sc_hd__buf_1 _4306_ (.A(_1772_),
    .X(_1773_));
 sky130_fd_sc_hd__buf_1 _4307_ (.A(_1039_),
    .X(_1774_));
 sky130_fd_sc_hd__inv_2 _4308_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][5] ),
    .Y(_1775_));
 sky130_fd_sc_hd__inv_2 _4309_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][1] ),
    .Y(_1776_));
 sky130_fd_sc_hd__buf_1 _4310_ (.A(_1041_),
    .X(_1777_));
 sky130_fd_sc_hd__inv_2 _4311_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][2] ),
    .Y(_1778_));
 sky130_fd_sc_hd__buf_1 _4312_ (.A(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__buf_1 _4313_ (.A(_1774_),
    .X(_1780_));
 sky130_fd_sc_hd__buf_1 _4314_ (.A(_1780_),
    .X(_1781_));
 sky130_fd_sc_hd__inv_2 _4315_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][6] ),
    .Y(_1782_));
 sky130_fd_sc_hd__buf_1 _4316_ (.A(_1035_),
    .X(_1783_));
 sky130_fd_sc_hd__buf_1 _4317_ (.A(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__buf_1 _4318_ (.A(_1048_),
    .X(_1785_));
 sky130_fd_sc_hd__buf_1 _4319_ (.A(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__buf_1 _4320_ (.A(_1770_),
    .X(_1787_));
 sky130_fd_sc_hd__buf_1 _4321_ (.A(_1787_),
    .X(_1788_));
 sky130_fd_sc_hd__nand2_2 _4322_ (.A(_1773_),
    .B(_1046_),
    .Y(_1789_));
 sky130_fd_sc_hd__buf_1 _4323_ (.A(_1777_),
    .X(_1790_));
 sky130_fd_sc_hd__buf_1 _4324_ (.A(_1776_),
    .X(_1791_));
 sky130_fd_sc_hd__nor2_2 _4325_ (.A(_1768_),
    .B(_1789_),
    .Y(_1792_));
 sky130_fd_sc_hd__buf_1 _4326_ (.A(_1049_),
    .X(_1793_));
 sky130_fd_sc_hd__buf_1 _4327_ (.A(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__buf_1 _4328_ (.A(_1794_),
    .X(_1795_));
 sky130_fd_sc_hd__nor2_2 _4329_ (.A(_1775_),
    .B(_1782_),
    .Y(_1796_));
 sky130_fd_sc_hd__buf_1 _4330_ (.A(_1771_),
    .X(_1797_));
 sky130_fd_sc_hd__and3_2 _4331_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][7] ),
    .B(_1796_),
    .C(_1792_),
    .X(_1798_));
 sky130_fd_sc_hd__buf_1 _4332_ (.A(_1798_),
    .X(_0218_));
 sky130_fd_sc_hd__buf_1 _4333_ (.A(_1795_),
    .X(_1799_));
 sky130_fd_sc_hd__buf_1 _4334_ (.A(_1786_),
    .X(_1800_));
 sky130_fd_sc_hd__or3b_2 _4335_ (.A(_0731_),
    .B(\tree_instances[18].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[18].u_tree.tree_state[0] ),
    .X(_1801_));
 sky130_fd_sc_hd__inv_2 _4336_ (.A(_1801_),
    .Y(_0022_));
 sky130_fd_sc_hd__and3b_2 _4337_ (.A_N(\tree_instances[20].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[20].u_tree.tree_state[0] ),
    .C(feature_valid),
    .X(_1802_));
 sky130_fd_sc_hd__buf_1 _4338_ (.A(_1802_),
    .X(_0028_));
 sky130_fd_sc_hd__buf_1 _4339_ (.A(_0730_),
    .X(_1803_));
 sky130_fd_sc_hd__or3b_2 _4340_ (.A(_1803_),
    .B(\tree_instances[2].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[2].u_tree.tree_state[0] ),
    .X(_1804_));
 sky130_fd_sc_hd__inv_2 _4341_ (.A(_1804_),
    .Y(_0030_));
 sky130_fd_sc_hd__and3b_2 _4342_ (.A_N(\tree_instances[17].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[17].u_tree.tree_state[0] ),
    .C(feature_valid),
    .X(_1805_));
 sky130_fd_sc_hd__buf_1 _4343_ (.A(_1805_),
    .X(_0020_));
 sky130_fd_sc_hd__and3b_2 _4344_ (.A_N(\tree_instances[3].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[3].u_tree.tree_state[0] ),
    .C(feature_valid),
    .X(_1806_));
 sky130_fd_sc_hd__buf_1 _4345_ (.A(_1806_),
    .X(_0032_));
 sky130_fd_sc_hd__or3b_2 _4346_ (.A(_1803_),
    .B(\tree_instances[4].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[4].u_tree.tree_state[0] ),
    .X(_1807_));
 sky130_fd_sc_hd__inv_2 _4347_ (.A(_1807_),
    .Y(_0034_));
 sky130_fd_sc_hd__or3b_2 _4348_ (.A(_1803_),
    .B(\tree_instances[5].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[5].u_tree.tree_state[0] ),
    .X(_1808_));
 sky130_fd_sc_hd__inv_2 _4349_ (.A(_1808_),
    .Y(_0036_));
 sky130_fd_sc_hd__or3b_2 _4350_ (.A(_1803_),
    .B(\tree_instances[16].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[16].u_tree.tree_state[0] ),
    .X(_1809_));
 sky130_fd_sc_hd__inv_2 _4351_ (.A(_1809_),
    .Y(_0018_));
 sky130_fd_sc_hd__or3b_2 _4352_ (.A(_1803_),
    .B(\tree_instances[12].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[12].u_tree.tree_state[0] ),
    .X(_1810_));
 sky130_fd_sc_hd__inv_2 _4353_ (.A(_1810_),
    .Y(_0010_));
 sky130_fd_sc_hd__or3b_2 _4354_ (.A(_1803_),
    .B(\tree_instances[6].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[6].u_tree.tree_state[0] ),
    .X(_1811_));
 sky130_fd_sc_hd__inv_2 _4355_ (.A(_1811_),
    .Y(_0038_));
 sky130_fd_sc_hd__or3b_2 _4356_ (.A(_1803_),
    .B(\tree_instances[7].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[7].u_tree.tree_state[0] ),
    .X(_1812_));
 sky130_fd_sc_hd__inv_2 _4357_ (.A(_1812_),
    .Y(_0040_));
 sky130_fd_sc_hd__or3b_2 _4358_ (.A(_1803_),
    .B(\tree_instances[8].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[8].u_tree.tree_state[0] ),
    .X(_1813_));
 sky130_fd_sc_hd__inv_2 _4359_ (.A(_1813_),
    .Y(_0042_));
 sky130_fd_sc_hd__or3b_2 _4360_ (.A(_1112_),
    .B(\tree_instances[9].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[9].u_tree.tree_state[0] ),
    .X(_1814_));
 sky130_fd_sc_hd__inv_2 _4361_ (.A(_1814_),
    .Y(_0044_));
 sky130_fd_sc_hd__and3b_2 _4362_ (.A_N(\tree_instances[15].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[15].u_tree.tree_state[0] ),
    .C(feature_valid),
    .X(_1815_));
 sky130_fd_sc_hd__buf_1 _4363_ (.A(_1815_),
    .X(_0016_));
 sky130_fd_sc_hd__or3b_2 _4364_ (.A(_1112_),
    .B(\tree_instances[11].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[11].u_tree.tree_state[0] ),
    .X(_1816_));
 sky130_fd_sc_hd__inv_2 _4365_ (.A(_1816_),
    .Y(_0008_));
 sky130_fd_sc_hd__or3b_2 _4366_ (.A(_1112_),
    .B(\tree_instances[14].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[14].u_tree.tree_state[0] ),
    .X(_1817_));
 sky130_fd_sc_hd__inv_2 _4367_ (.A(_1817_),
    .Y(_0014_));
 sky130_fd_sc_hd__or3b_2 _4368_ (.A(_1112_),
    .B(\tree_instances[0].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[0].u_tree.tree_state[0] ),
    .X(_1818_));
 sky130_fd_sc_hd__inv_2 _4369_ (.A(_1818_),
    .Y(_0004_));
 sky130_fd_sc_hd__or3b_2 _4370_ (.A(_1112_),
    .B(\tree_instances[10].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[10].u_tree.tree_state[0] ),
    .X(_1819_));
 sky130_fd_sc_hd__inv_2 _4371_ (.A(_1819_),
    .Y(_0006_));
 sky130_fd_sc_hd__or3b_2 _4372_ (.A(_1112_),
    .B(\tree_instances[1].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[1].u_tree.tree_state[0] ),
    .X(_1820_));
 sky130_fd_sc_hd__inv_2 _4373_ (.A(_1820_),
    .Y(_0026_));
 sky130_fd_sc_hd__inv_2 _4374_ (.A(_0865_),
    .Y(_1821_));
 sky130_fd_sc_hd__nor2_2 _4375_ (.A(_1821_),
    .B(_0883_),
    .Y(_0025_));
 sky130_fd_sc_hd__inv_2 _4376_ (.A(\tree_instances[13].u_tree.tree_state[0] ),
    .Y(_1822_));
 sky130_fd_sc_hd__or2_2 _4377_ (.A(_1822_),
    .B(_1113_),
    .X(_1823_));
 sky130_fd_sc_hd__buf_1 _4378_ (.A(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__inv_2 _4379_ (.A(_1824_),
    .Y(_0012_));
 sky130_fd_sc_hd__or3b_2 _4380_ (.A(_1112_),
    .B(\tree_instances[19].u_tree.pipeline_valid[0] ),
    .C_N(\tree_instances[19].u_tree.tree_state[0] ),
    .X(_1825_));
 sky130_fd_sc_hd__inv_2 _4381_ (.A(_1825_),
    .Y(_0024_));
 sky130_fd_sc_hd__buf_1 _4382_ (.A(\tree_instances[0].u_tree.frame_id_in[0] ),
    .X(_1826_));
 sky130_fd_sc_hd__buf_1 _4383_ (.A(_1826_),
    .X(_1827_));
 sky130_fd_sc_hd__mux2_2 _4384_ (.A0(\tree_instances[7].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1827_),
    .S(_0040_),
    .X(_1828_));
 sky130_fd_sc_hd__buf_1 _4385_ (.A(_1828_),
    .X(_0108_));
 sky130_fd_sc_hd__buf_1 _4386_ (.A(\tree_instances[0].u_tree.frame_id_in[1] ),
    .X(_1829_));
 sky130_fd_sc_hd__buf_1 _4387_ (.A(_1829_),
    .X(_1830_));
 sky130_fd_sc_hd__mux2_2 _4388_ (.A0(\tree_instances[7].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1830_),
    .S(_0040_),
    .X(_1831_));
 sky130_fd_sc_hd__buf_1 _4389_ (.A(_1831_),
    .X(_0109_));
 sky130_fd_sc_hd__buf_1 _4390_ (.A(\tree_instances[0].u_tree.frame_id_in[2] ),
    .X(_1832_));
 sky130_fd_sc_hd__mux2_2 _4391_ (.A0(\tree_instances[7].u_tree.pipeline_frame_id[0][2] ),
    .A1(_1832_),
    .S(_0040_),
    .X(_1833_));
 sky130_fd_sc_hd__buf_1 _4392_ (.A(_1833_),
    .X(_0110_));
 sky130_fd_sc_hd__buf_1 _4393_ (.A(\tree_instances[0].u_tree.frame_id_in[3] ),
    .X(_1834_));
 sky130_fd_sc_hd__buf_1 _4394_ (.A(_1834_),
    .X(_1835_));
 sky130_fd_sc_hd__mux2_2 _4395_ (.A0(\tree_instances[7].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1835_),
    .S(_0040_),
    .X(_1836_));
 sky130_fd_sc_hd__buf_1 _4396_ (.A(_1836_),
    .X(_0111_));
 sky130_fd_sc_hd__buf_1 _4397_ (.A(\tree_instances[0].u_tree.frame_id_in[4] ),
    .X(_1837_));
 sky130_fd_sc_hd__mux2_2 _4398_ (.A0(\tree_instances[7].u_tree.pipeline_frame_id[0][4] ),
    .A1(_1837_),
    .S(_0040_),
    .X(_1838_));
 sky130_fd_sc_hd__buf_1 _4399_ (.A(_1838_),
    .X(_0112_));
 sky130_fd_sc_hd__or3_2 _4400_ (.A(\tree_instances[7].u_tree.tree_state[2] ),
    .B(\tree_instances[7].u_tree.tree_state[1] ),
    .C(_1812_),
    .X(_1839_));
 sky130_fd_sc_hd__buf_1 _4401_ (.A(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__mux2_2 _4402_ (.A0(\tree_instances[7].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[7].u_tree.pipeline_frame_id[0][0] ),
    .S(_0970_),
    .X(_1841_));
 sky130_fd_sc_hd__buf_1 _4403_ (.A(_1841_),
    .X(_0113_));
 sky130_fd_sc_hd__mux2_2 _4404_ (.A0(\tree_instances[7].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[7].u_tree.pipeline_frame_id[0][1] ),
    .S(_0970_),
    .X(_1842_));
 sky130_fd_sc_hd__buf_1 _4405_ (.A(_1842_),
    .X(_0114_));
 sky130_fd_sc_hd__mux2_2 _4406_ (.A0(\tree_instances[7].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[7].u_tree.pipeline_frame_id[0][2] ),
    .S(_0970_),
    .X(_1843_));
 sky130_fd_sc_hd__buf_1 _4407_ (.A(_1843_),
    .X(_0115_));
 sky130_fd_sc_hd__mux2_2 _4408_ (.A0(\tree_instances[7].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[7].u_tree.pipeline_frame_id[0][3] ),
    .S(_0970_),
    .X(_1844_));
 sky130_fd_sc_hd__buf_1 _4409_ (.A(_1844_),
    .X(_0116_));
 sky130_fd_sc_hd__mux2_2 _4410_ (.A0(\tree_instances[7].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[7].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[7].u_tree.tree_state[3] ),
    .X(_1845_));
 sky130_fd_sc_hd__buf_1 _4411_ (.A(_1845_),
    .X(_0117_));
 sky130_fd_sc_hd__buf_1 _4412_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][0] ),
    .X(_1846_));
 sky130_fd_sc_hd__buf_1 _4413_ (.A(_1846_),
    .X(_1847_));
 sky130_fd_sc_hd__buf_1 _4414_ (.A(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__buf_1 _4415_ (.A(_1848_),
    .X(_1849_));
 sky130_fd_sc_hd__or3_2 _4416_ (.A(\tree_instances[6].u_tree.tree_state[1] ),
    .B(\tree_instances[6].u_tree.tree_state[2] ),
    .C(_1811_),
    .X(_1850_));
 sky130_fd_sc_hd__buf_1 _4417_ (.A(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__and2_2 _4418_ (.A(_1849_),
    .B(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__buf_1 _4419_ (.A(_1852_),
    .X(_0118_));
 sky130_fd_sc_hd__buf_1 _4420_ (.A(_0977_),
    .X(_1853_));
 sky130_fd_sc_hd__buf_1 _4421_ (.A(_1853_),
    .X(_1854_));
 sky130_fd_sc_hd__buf_1 _4422_ (.A(_1854_),
    .X(_1855_));
 sky130_fd_sc_hd__buf_1 _4423_ (.A(_1855_),
    .X(_1856_));
 sky130_fd_sc_hd__and2_2 _4424_ (.A(_1856_),
    .B(_1851_),
    .X(_1857_));
 sky130_fd_sc_hd__buf_1 _4425_ (.A(_1857_),
    .X(_0119_));
 sky130_fd_sc_hd__buf_1 _4426_ (.A(_0985_),
    .X(_1858_));
 sky130_fd_sc_hd__and2_2 _4427_ (.A(_1858_),
    .B(_1851_),
    .X(_1859_));
 sky130_fd_sc_hd__buf_1 _4428_ (.A(_1859_),
    .X(_0120_));
 sky130_fd_sc_hd__buf_1 _4429_ (.A(_0981_),
    .X(_1860_));
 sky130_fd_sc_hd__buf_1 _4430_ (.A(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__buf_1 _4431_ (.A(_1861_),
    .X(_1862_));
 sky130_fd_sc_hd__buf_1 _4432_ (.A(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__and2_2 _4433_ (.A(_1863_),
    .B(_1851_),
    .X(_1864_));
 sky130_fd_sc_hd__buf_1 _4434_ (.A(_1864_),
    .X(_0121_));
 sky130_fd_sc_hd__buf_1 _4435_ (.A(_0973_),
    .X(_1865_));
 sky130_fd_sc_hd__buf_1 _4436_ (.A(_1865_),
    .X(_1866_));
 sky130_fd_sc_hd__buf_1 _4437_ (.A(_1866_),
    .X(_1867_));
 sky130_fd_sc_hd__buf_1 _4438_ (.A(_1867_),
    .X(_1868_));
 sky130_fd_sc_hd__and2_2 _4439_ (.A(_1868_),
    .B(_1851_),
    .X(_1869_));
 sky130_fd_sc_hd__buf_1 _4440_ (.A(_1869_),
    .X(_0122_));
 sky130_fd_sc_hd__buf_1 _4441_ (.A(_0972_),
    .X(_1870_));
 sky130_fd_sc_hd__buf_1 _4442_ (.A(_1870_),
    .X(_1871_));
 sky130_fd_sc_hd__buf_1 _4443_ (.A(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__and2_2 _4444_ (.A(_1872_),
    .B(_1851_),
    .X(_1873_));
 sky130_fd_sc_hd__buf_1 _4445_ (.A(_1873_),
    .X(_0123_));
 sky130_fd_sc_hd__buf_1 _4446_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][6] ),
    .X(_1874_));
 sky130_fd_sc_hd__buf_1 _4447_ (.A(_1874_),
    .X(_1875_));
 sky130_fd_sc_hd__buf_1 _4448_ (.A(_1875_),
    .X(_1876_));
 sky130_fd_sc_hd__buf_1 _4449_ (.A(_1876_),
    .X(_1877_));
 sky130_fd_sc_hd__and2_2 _4450_ (.A(_1877_),
    .B(_1851_),
    .X(_1878_));
 sky130_fd_sc_hd__buf_1 _4451_ (.A(_1878_),
    .X(_0124_));
 sky130_fd_sc_hd__buf_1 _4452_ (.A(\tree_instances[6].u_tree.pipeline_current_node[0][7] ),
    .X(_1879_));
 sky130_fd_sc_hd__buf_1 _4453_ (.A(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__and2_2 _4454_ (.A(_1880_),
    .B(_1850_),
    .X(_1881_));
 sky130_fd_sc_hd__buf_1 _4455_ (.A(_1881_),
    .X(_0125_));
 sky130_fd_sc_hd__and2_2 _4456_ (.A(_1233_),
    .B(_1850_),
    .X(_1882_));
 sky130_fd_sc_hd__buf_1 _4457_ (.A(_1882_),
    .X(_0126_));
 sky130_fd_sc_hd__nand2_2 _4458_ (.A(\tree_instances[7].u_tree.tree_state[0] ),
    .B(_0969_),
    .Y(_1883_));
 sky130_fd_sc_hd__a22o_2 _4459_ (.A1(_0970_),
    .A2(_1883_),
    .B1(_1812_),
    .B2(\tree_instances[7].u_tree.ready_for_next ),
    .X(_0127_));
 sky130_fd_sc_hd__nand2_2 _4460_ (.A(\tree_instances[18].u_tree.tree_state[0] ),
    .B(_0752_),
    .Y(_1884_));
 sky130_fd_sc_hd__o2bb2a_2 _4461_ (.A1_N(_0753_),
    .A2_N(_1884_),
    .B1(_0022_),
    .B2(\tree_instances[18].u_tree.pipeline_valid[0] ),
    .X(_0128_));
 sky130_fd_sc_hd__buf_1 _4462_ (.A(_0713_),
    .X(_1885_));
 sky130_fd_sc_hd__buf_1 _4463_ (.A(_0716_),
    .X(_1886_));
 sky130_fd_sc_hd__buf_1 _4464_ (.A(_1886_),
    .X(_1887_));
 sky130_fd_sc_hd__buf_1 _4465_ (.A(_1887_),
    .X(_1888_));
 sky130_fd_sc_hd__buf_1 _4466_ (.A(_0724_),
    .X(_1889_));
 sky130_fd_sc_hd__buf_1 _4467_ (.A(_1889_),
    .X(_1890_));
 sky130_fd_sc_hd__buf_1 _4468_ (.A(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__buf_1 _4469_ (.A(_0715_),
    .X(_1892_));
 sky130_fd_sc_hd__buf_1 _4470_ (.A(_1892_),
    .X(_1893_));
 sky130_fd_sc_hd__buf_1 _4471_ (.A(_1893_),
    .X(_1894_));
 sky130_fd_sc_hd__buf_1 _4472_ (.A(\tree_instances[8].u_tree.tree_state[2] ),
    .X(_1895_));
 sky130_fd_sc_hd__a22o_2 _4473_ (.A1(\tree_instances[8].u_tree.tree_state[1] ),
    .A2(\tree_instances[8].u_tree.current_node_data[12] ),
    .B1(\tree_instances[8].u_tree.node_data[12] ),
    .B2(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__nand2_2 _4474_ (.A(\tree_instances[8].u_tree.tree_state[0] ),
    .B(_0999_),
    .Y(_1897_));
 sky130_fd_sc_hd__o31ai_2 _4475_ (.A1(\tree_instances[8].u_tree.tree_state[0] ),
    .A2(\tree_instances[8].u_tree.tree_state[2] ),
    .A3(\tree_instances[8].u_tree.tree_state[1] ),
    .B1(_1897_),
    .Y(_1898_));
 sky130_fd_sc_hd__nor2_2 _4476_ (.A(_0041_),
    .B(_1898_),
    .Y(_1899_));
 sky130_fd_sc_hd__mux2_2 _4477_ (.A0(\tree_instances[8].u_tree.pipeline_prediction[0][0] ),
    .A1(_1896_),
    .S(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__buf_1 _4478_ (.A(_1900_),
    .X(_0129_));
 sky130_fd_sc_hd__buf_1 _4479_ (.A(\tree_instances[8].u_tree.read_enable ),
    .X(_1901_));
 sky130_fd_sc_hd__buf_1 _4480_ (.A(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__nand2_2 _4481_ (.A(_1770_),
    .B(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .Y(_1903_));
 sky130_fd_sc_hd__or2_2 _4482_ (.A(_1765_),
    .B(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .X(_1904_));
 sky130_fd_sc_hd__nand2_2 _4483_ (.A(_1046_),
    .B(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .Y(_1905_));
 sky130_fd_sc_hd__or2_2 _4484_ (.A(_1046_),
    .B(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .X(_1906_));
 sky130_fd_sc_hd__xor2_2 _4485_ (.A(\tree_instances[8].u_tree.pipeline_current_node[0][7] ),
    .B(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .X(_1907_));
 sky130_fd_sc_hd__a221o_2 _4486_ (.A1(_1903_),
    .A2(_1904_),
    .B1(_1905_),
    .B2(_1906_),
    .C1(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__inv_2 _4487_ (.A(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .Y(_1909_));
 sky130_fd_sc_hd__inv_2 _4488_ (.A(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .Y(_1910_));
 sky130_fd_sc_hd__o22a_2 _4489_ (.A1(_1791_),
    .A2(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .B1(_1910_),
    .B2(_1036_),
    .X(_1911_));
 sky130_fd_sc_hd__o21ai_2 _4490_ (.A1(_1774_),
    .A2(_1909_),
    .B1(_1911_),
    .Y(_1912_));
 sky130_fd_sc_hd__a2bb2o_2 _4491_ (.A1_N(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .A2_N(_1778_),
    .B1(_1774_),
    .B2(_1909_),
    .X(_1913_));
 sky130_fd_sc_hd__a221o_2 _4492_ (.A1(_1779_),
    .A2(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .B1(_1910_),
    .B2(_1036_),
    .C1(_1913_),
    .X(_1914_));
 sky130_fd_sc_hd__o21ai_2 _4493_ (.A1(_1775_),
    .A2(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .B1(\tree_instances[8].u_tree.u_tree_weight_rom.cache_valid ),
    .Y(_1915_));
 sky130_fd_sc_hd__a221o_2 _4494_ (.A1(_1791_),
    .A2(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .B1(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .B2(_1775_),
    .C1(_1915_),
    .X(_1916_));
 sky130_fd_sc_hd__or4_2 _4495_ (.A(_1908_),
    .B(_1912_),
    .C(_1914_),
    .D(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__buf_1 _4496_ (.A(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__a21o_2 _4497_ (.A1(_1902_),
    .A2(_1918_),
    .B1(\tree_instances[8].u_tree.u_tree_weight_rom.cache_valid ),
    .X(_0130_));
 sky130_fd_sc_hd__and2_2 _4498_ (.A(_1290_),
    .B(_1840_),
    .X(_1919_));
 sky130_fd_sc_hd__buf_1 _4499_ (.A(_1919_),
    .X(_0131_));
 sky130_fd_sc_hd__and2_2 _4500_ (.A(_1304_),
    .B(_1840_),
    .X(_1920_));
 sky130_fd_sc_hd__buf_1 _4501_ (.A(_1920_),
    .X(_0132_));
 sky130_fd_sc_hd__and2_2 _4502_ (.A(_1310_),
    .B(_1840_),
    .X(_1921_));
 sky130_fd_sc_hd__buf_1 _4503_ (.A(_1921_),
    .X(_0133_));
 sky130_fd_sc_hd__and2_2 _4504_ (.A(_1309_),
    .B(_1840_),
    .X(_1922_));
 sky130_fd_sc_hd__buf_1 _4505_ (.A(_1922_),
    .X(_0134_));
 sky130_fd_sc_hd__and2_2 _4506_ (.A(_1305_),
    .B(_1840_),
    .X(_1923_));
 sky130_fd_sc_hd__buf_1 _4507_ (.A(_1923_),
    .X(_0135_));
 sky130_fd_sc_hd__and2_2 _4508_ (.A(_1300_),
    .B(_1840_),
    .X(_1924_));
 sky130_fd_sc_hd__buf_1 _4509_ (.A(_1924_),
    .X(_0136_));
 sky130_fd_sc_hd__and2_2 _4510_ (.A(_1313_),
    .B(_1840_),
    .X(_1925_));
 sky130_fd_sc_hd__buf_1 _4511_ (.A(_1925_),
    .X(_0137_));
 sky130_fd_sc_hd__and2_2 _4512_ (.A(_1302_),
    .B(_1839_),
    .X(_1926_));
 sky130_fd_sc_hd__buf_1 _4513_ (.A(_1926_),
    .X(_0138_));
 sky130_fd_sc_hd__mux2_2 _4514_ (.A0(\tree_instances[8].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1827_),
    .S(_0042_),
    .X(_1927_));
 sky130_fd_sc_hd__buf_1 _4515_ (.A(_1927_),
    .X(_0139_));
 sky130_fd_sc_hd__mux2_2 _4516_ (.A0(\tree_instances[8].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1830_),
    .S(_0042_),
    .X(_1928_));
 sky130_fd_sc_hd__buf_1 _4517_ (.A(_1928_),
    .X(_0140_));
 sky130_fd_sc_hd__mux2_2 _4518_ (.A0(\tree_instances[8].u_tree.pipeline_frame_id[0][2] ),
    .A1(_1832_),
    .S(_0042_),
    .X(_1929_));
 sky130_fd_sc_hd__buf_1 _4519_ (.A(_1929_),
    .X(_0141_));
 sky130_fd_sc_hd__mux2_2 _4520_ (.A0(\tree_instances[8].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1835_),
    .S(_0042_),
    .X(_1930_));
 sky130_fd_sc_hd__buf_1 _4521_ (.A(_1930_),
    .X(_0142_));
 sky130_fd_sc_hd__mux2_2 _4522_ (.A0(\tree_instances[8].u_tree.pipeline_frame_id[0][4] ),
    .A1(_1837_),
    .S(_0042_),
    .X(_1931_));
 sky130_fd_sc_hd__buf_1 _4523_ (.A(_1931_),
    .X(_0143_));
 sky130_fd_sc_hd__inv_2 _4524_ (.A(\tree_instances[8].u_tree.read_enable ),
    .Y(_1932_));
 sky130_fd_sc_hd__buf_1 _4525_ (.A(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__buf_1 _4526_ (.A(_1933_),
    .X(_1934_));
 sky130_fd_sc_hd__o21ba_2 _4527_ (.A1(\tree_instances[8].u_tree.tree_state[0] ),
    .A2(_1034_),
    .B1_N(\tree_instances[8].u_tree.tree_state[1] ),
    .X(_1935_));
 sky130_fd_sc_hd__or3_2 _4528_ (.A(\tree_instances[8].u_tree.tree_state[2] ),
    .B(\tree_instances[8].u_tree.tree_state[1] ),
    .C(_1813_),
    .X(_1936_));
 sky130_fd_sc_hd__buf_1 _4529_ (.A(_1936_),
    .X(_1937_));
 sky130_fd_sc_hd__o21ai_2 _4530_ (.A1(_1934_),
    .A2(_1935_),
    .B1(_1937_),
    .Y(_0144_));
 sky130_fd_sc_hd__mux2_2 _4531_ (.A0(\tree_instances[8].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[8].u_tree.pipeline_frame_id[0][0] ),
    .S(_1000_),
    .X(_1938_));
 sky130_fd_sc_hd__buf_1 _4532_ (.A(_1938_),
    .X(_0145_));
 sky130_fd_sc_hd__mux2_2 _4533_ (.A0(\tree_instances[8].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[8].u_tree.pipeline_frame_id[0][1] ),
    .S(_1000_),
    .X(_1939_));
 sky130_fd_sc_hd__buf_1 _4534_ (.A(_1939_),
    .X(_0146_));
 sky130_fd_sc_hd__mux2_2 _4535_ (.A0(\tree_instances[8].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[8].u_tree.pipeline_frame_id[0][2] ),
    .S(_1000_),
    .X(_1940_));
 sky130_fd_sc_hd__buf_1 _4536_ (.A(_1940_),
    .X(_0147_));
 sky130_fd_sc_hd__mux2_2 _4537_ (.A0(\tree_instances[8].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[8].u_tree.pipeline_frame_id[0][3] ),
    .S(_1000_),
    .X(_1941_));
 sky130_fd_sc_hd__buf_1 _4538_ (.A(_1941_),
    .X(_0148_));
 sky130_fd_sc_hd__mux2_2 _4539_ (.A0(\tree_instances[8].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[8].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[8].u_tree.tree_state[3] ),
    .X(_1942_));
 sky130_fd_sc_hd__buf_1 _4540_ (.A(_1942_),
    .X(_0149_));
 sky130_fd_sc_hd__mux2_2 _4541_ (.A0(\tree_instances[8].u_tree.prediction_out ),
    .A1(\tree_instances[8].u_tree.pipeline_prediction[0][0] ),
    .S(\tree_instances[8].u_tree.tree_state[3] ),
    .X(_1943_));
 sky130_fd_sc_hd__buf_1 _4542_ (.A(_1943_),
    .X(_0150_));
 sky130_fd_sc_hd__a22o_2 _4543_ (.A1(_1000_),
    .A2(_1897_),
    .B1(_1813_),
    .B2(\tree_instances[8].u_tree.ready_for_next ),
    .X(_0151_));
 sky130_fd_sc_hd__or3_2 _4544_ (.A(\tree_instances[9].u_tree.tree_state[1] ),
    .B(\tree_instances[9].u_tree.tree_state[2] ),
    .C(_1814_),
    .X(_1944_));
 sky130_fd_sc_hd__buf_1 _4545_ (.A(_1944_),
    .X(_1945_));
 sky130_fd_sc_hd__and2_2 _4546_ (.A(_1750_),
    .B(_1945_),
    .X(_1946_));
 sky130_fd_sc_hd__buf_1 _4547_ (.A(_1946_),
    .X(_0152_));
 sky130_fd_sc_hd__and2_2 _4548_ (.A(_1742_),
    .B(_1945_),
    .X(_1947_));
 sky130_fd_sc_hd__buf_1 _4549_ (.A(_1947_),
    .X(_0153_));
 sky130_fd_sc_hd__and2_2 _4550_ (.A(_1760_),
    .B(_1945_),
    .X(_1948_));
 sky130_fd_sc_hd__buf_1 _4551_ (.A(_1948_),
    .X(_0154_));
 sky130_fd_sc_hd__and2_2 _4552_ (.A(_1757_),
    .B(_1945_),
    .X(_1949_));
 sky130_fd_sc_hd__buf_1 _4553_ (.A(_1949_),
    .X(_0155_));
 sky130_fd_sc_hd__and2_2 _4554_ (.A(_1759_),
    .B(_1945_),
    .X(_1950_));
 sky130_fd_sc_hd__buf_1 _4555_ (.A(_1950_),
    .X(_0156_));
 sky130_fd_sc_hd__and2_2 _4556_ (.A(_1749_),
    .B(_1945_),
    .X(_1951_));
 sky130_fd_sc_hd__buf_1 _4557_ (.A(_1951_),
    .X(_0157_));
 sky130_fd_sc_hd__and2_2 _4558_ (.A(_1755_),
    .B(_1945_),
    .X(_1952_));
 sky130_fd_sc_hd__buf_1 _4559_ (.A(_1952_),
    .X(_0158_));
 sky130_fd_sc_hd__and2_2 _4560_ (.A(_1752_),
    .B(_1944_),
    .X(_1953_));
 sky130_fd_sc_hd__buf_1 _4561_ (.A(_1953_),
    .X(_0159_));
 sky130_fd_sc_hd__o2bb2a_2 _4562_ (.A1_N(_1197_),
    .A2_N(_1198_),
    .B1(_0028_),
    .B2(\tree_instances[20].u_tree.pipeline_valid[0] ),
    .X(_0160_));
 sky130_fd_sc_hd__and4_2 _4563_ (.A(_1724_),
    .B(_1701_),
    .C(_1706_),
    .D(_1722_),
    .X(_1954_));
 sky130_fd_sc_hd__buf_1 _4564_ (.A(_1954_),
    .X(_0161_));
 sky130_fd_sc_hd__nand2_2 _4565_ (.A(\tree_instances[4].u_tree.tree_state[0] ),
    .B(_0848_),
    .Y(_1955_));
 sky130_fd_sc_hd__o2bb2a_2 _4566_ (.A1_N(_0849_),
    .A2_N(_1955_),
    .B1(_0034_),
    .B2(\tree_instances[4].u_tree.pipeline_valid[0] ),
    .X(_0162_));
 sky130_fd_sc_hd__nand2_2 _4567_ (.A(\tree_instances[8].u_tree.read_enable ),
    .B(_1917_),
    .Y(_1956_));
 sky130_fd_sc_hd__buf_1 _4568_ (.A(_1956_),
    .X(_1957_));
 sky130_fd_sc_hd__mux2_2 _4569_ (.A0(_1781_),
    .A1(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .S(_1957_),
    .X(_1958_));
 sky130_fd_sc_hd__buf_1 _4570_ (.A(_1958_),
    .X(_0163_));
 sky130_fd_sc_hd__mux2_2 _4571_ (.A0(_1790_),
    .A1(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .S(_1956_),
    .X(_1959_));
 sky130_fd_sc_hd__buf_1 _4572_ (.A(_1959_),
    .X(_0164_));
 sky130_fd_sc_hd__mux2_2 _4573_ (.A0(_1797_),
    .A1(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .S(_1956_),
    .X(_1960_));
 sky130_fd_sc_hd__buf_1 _4574_ (.A(_1960_),
    .X(_0165_));
 sky130_fd_sc_hd__mux2_2 _4575_ (.A0(_1788_),
    .A1(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .S(_1956_),
    .X(_1961_));
 sky130_fd_sc_hd__buf_1 _4576_ (.A(_1961_),
    .X(_0166_));
 sky130_fd_sc_hd__mux2_2 _4577_ (.A0(_1800_),
    .A1(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .S(_1956_),
    .X(_1962_));
 sky130_fd_sc_hd__buf_1 _4578_ (.A(_1962_),
    .X(_0167_));
 sky130_fd_sc_hd__mux2_2 _4579_ (.A0(_1799_),
    .A1(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .S(_1956_),
    .X(_1963_));
 sky130_fd_sc_hd__buf_1 _4580_ (.A(_1963_),
    .X(_0168_));
 sky130_fd_sc_hd__mux2_2 _4581_ (.A0(_1764_),
    .A1(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .S(_1956_),
    .X(_1964_));
 sky130_fd_sc_hd__buf_1 _4582_ (.A(_1964_),
    .X(_0169_));
 sky130_fd_sc_hd__mux2_2 _4583_ (.A0(_1784_),
    .A1(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .S(_1956_),
    .X(_1965_));
 sky130_fd_sc_hd__buf_1 _4584_ (.A(_1965_),
    .X(_0170_));
 sky130_fd_sc_hd__buf_1 _4585_ (.A(_1957_),
    .X(_1966_));
 sky130_fd_sc_hd__and3_2 _4586_ (.A(_1902_),
    .B(\tree_instances[8].u_tree.u_tree_weight_rom.gen_tree_8.u_tree_rom.node_data[12] ),
    .C(_1918_),
    .X(_1967_));
 sky130_fd_sc_hd__a21o_2 _4587_ (.A1(\tree_instances[8].u_tree.u_tree_weight_rom.cached_data[12] ),
    .A2(_1966_),
    .B1(_1967_),
    .X(_0171_));
 sky130_fd_sc_hd__buf_1 _4588_ (.A(_1917_),
    .X(_1968_));
 sky130_fd_sc_hd__mux2_2 _4589_ (.A0(\tree_instances[9].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1827_),
    .S(_0044_),
    .X(_1969_));
 sky130_fd_sc_hd__buf_1 _4590_ (.A(_1969_),
    .X(_0172_));
 sky130_fd_sc_hd__mux2_2 _4591_ (.A0(\tree_instances[9].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1830_),
    .S(_0044_),
    .X(_1970_));
 sky130_fd_sc_hd__buf_1 _4592_ (.A(_1970_),
    .X(_0173_));
 sky130_fd_sc_hd__mux2_2 _4593_ (.A0(\tree_instances[9].u_tree.pipeline_frame_id[0][2] ),
    .A1(_1832_),
    .S(_0044_),
    .X(_1971_));
 sky130_fd_sc_hd__buf_1 _4594_ (.A(_1971_),
    .X(_0174_));
 sky130_fd_sc_hd__mux2_2 _4595_ (.A0(\tree_instances[9].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1835_),
    .S(_0044_),
    .X(_1972_));
 sky130_fd_sc_hd__buf_1 _4596_ (.A(_1972_),
    .X(_0175_));
 sky130_fd_sc_hd__mux2_2 _4597_ (.A0(\tree_instances[9].u_tree.pipeline_frame_id[0][4] ),
    .A1(_1837_),
    .S(_0044_),
    .X(_1973_));
 sky130_fd_sc_hd__buf_1 _4598_ (.A(_1973_),
    .X(_0176_));
 sky130_fd_sc_hd__mux2_2 _4599_ (.A0(\tree_instances[8].u_tree.current_node_data[12] ),
    .A1(\tree_instances[8].u_tree.node_data[12] ),
    .S(_1034_),
    .X(_1974_));
 sky130_fd_sc_hd__buf_1 _4600_ (.A(_1974_),
    .X(_0177_));
 sky130_fd_sc_hd__mux2_2 _4601_ (.A0(\tree_instances[9].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[9].u_tree.pipeline_frame_id[0][0] ),
    .S(_1025_),
    .X(_1975_));
 sky130_fd_sc_hd__buf_1 _4602_ (.A(_1975_),
    .X(_0178_));
 sky130_fd_sc_hd__mux2_2 _4603_ (.A0(\tree_instances[9].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[9].u_tree.pipeline_frame_id[0][1] ),
    .S(_1025_),
    .X(_1976_));
 sky130_fd_sc_hd__buf_1 _4604_ (.A(_1976_),
    .X(_0179_));
 sky130_fd_sc_hd__mux2_2 _4605_ (.A0(\tree_instances[9].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[9].u_tree.pipeline_frame_id[0][2] ),
    .S(_1025_),
    .X(_1977_));
 sky130_fd_sc_hd__buf_1 _4606_ (.A(_1977_),
    .X(_0180_));
 sky130_fd_sc_hd__mux2_2 _4607_ (.A0(\tree_instances[9].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[9].u_tree.pipeline_frame_id[0][3] ),
    .S(_1025_),
    .X(_1978_));
 sky130_fd_sc_hd__buf_1 _4608_ (.A(_1978_),
    .X(_0181_));
 sky130_fd_sc_hd__mux2_2 _4609_ (.A0(\tree_instances[9].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[9].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[9].u_tree.tree_state[3] ),
    .X(_1979_));
 sky130_fd_sc_hd__buf_1 _4610_ (.A(_1979_),
    .X(_0182_));
 sky130_fd_sc_hd__and2_2 _4611_ (.A(_1781_),
    .B(_1937_),
    .X(_1980_));
 sky130_fd_sc_hd__buf_1 _4612_ (.A(_1980_),
    .X(_0183_));
 sky130_fd_sc_hd__and2_2 _4613_ (.A(_1790_),
    .B(_1937_),
    .X(_1981_));
 sky130_fd_sc_hd__buf_1 _4614_ (.A(_1981_),
    .X(_0184_));
 sky130_fd_sc_hd__and2_2 _4615_ (.A(_1797_),
    .B(_1937_),
    .X(_1982_));
 sky130_fd_sc_hd__buf_1 _4616_ (.A(_1982_),
    .X(_0185_));
 sky130_fd_sc_hd__and2_2 _4617_ (.A(_1788_),
    .B(_1937_),
    .X(_1983_));
 sky130_fd_sc_hd__buf_1 _4618_ (.A(_1983_),
    .X(_0186_));
 sky130_fd_sc_hd__and2_2 _4619_ (.A(_1800_),
    .B(_1937_),
    .X(_1984_));
 sky130_fd_sc_hd__buf_1 _4620_ (.A(_1984_),
    .X(_0187_));
 sky130_fd_sc_hd__and2_2 _4621_ (.A(_1799_),
    .B(_1937_),
    .X(_1985_));
 sky130_fd_sc_hd__buf_1 _4622_ (.A(_1985_),
    .X(_0188_));
 sky130_fd_sc_hd__and2_2 _4623_ (.A(_1764_),
    .B(_1937_),
    .X(_1986_));
 sky130_fd_sc_hd__buf_1 _4624_ (.A(_1986_),
    .X(_0189_));
 sky130_fd_sc_hd__and2_2 _4625_ (.A(_1784_),
    .B(_1936_),
    .X(_1987_));
 sky130_fd_sc_hd__buf_1 _4626_ (.A(_1987_),
    .X(_0190_));
 sky130_fd_sc_hd__nand2_2 _4627_ (.A(\tree_instances[9].u_tree.tree_state[0] ),
    .B(_1024_),
    .Y(_1988_));
 sky130_fd_sc_hd__a22o_2 _4628_ (.A1(_1025_),
    .A2(_1988_),
    .B1(_1814_),
    .B2(\tree_instances[9].u_tree.ready_for_next ),
    .X(_0191_));
 sky130_fd_sc_hd__nand2_2 _4629_ (.A(\tree_instances[19].u_tree.tree_state[0] ),
    .B(_1251_),
    .Y(_1989_));
 sky130_fd_sc_hd__o2bb2a_2 _4630_ (.A1_N(_1252_),
    .A2_N(_1989_),
    .B1(_0024_),
    .B2(\tree_instances[19].u_tree.pipeline_valid[0] ),
    .X(_0192_));
 sky130_fd_sc_hd__a22o_2 _4631_ (.A1(\tree_instances[10].u_tree.tree_state[1] ),
    .A2(\tree_instances[10].u_tree.current_node_data[12] ),
    .B1(\tree_instances[10].u_tree.node_data[12] ),
    .B2(_1171_),
    .X(_1990_));
 sky130_fd_sc_hd__nand2_2 _4632_ (.A(\tree_instances[10].u_tree.tree_state[0] ),
    .B(_1135_),
    .Y(_1991_));
 sky130_fd_sc_hd__o311a_2 _4633_ (.A1(\tree_instances[10].u_tree.tree_state[0] ),
    .A2(\tree_instances[10].u_tree.tree_state[1] ),
    .A3(\tree_instances[10].u_tree.tree_state[2] ),
    .B1(_1991_),
    .C1(_1170_),
    .X(_1992_));
 sky130_fd_sc_hd__mux2_2 _4634_ (.A0(\tree_instances[10].u_tree.pipeline_prediction[0][0] ),
    .A1(_1990_),
    .S(_1992_),
    .X(_1993_));
 sky130_fd_sc_hd__buf_1 _4635_ (.A(_1993_),
    .X(_0193_));
 sky130_fd_sc_hd__inv_2 _4636_ (.A(\tree_instances[10].u_tree.u_tree_weight_rom.cache_valid ),
    .Y(_1994_));
 sky130_fd_sc_hd__inv_2 _4637_ (.A(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .Y(_1995_));
 sky130_fd_sc_hd__inv_2 _4638_ (.A(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .Y(_1996_));
 sky130_fd_sc_hd__xor2_2 _4639_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][5] ),
    .B(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .X(_1997_));
 sky130_fd_sc_hd__a221o_2 _4640_ (.A1(_1597_),
    .A2(_1995_),
    .B1(_1996_),
    .B2(\tree_instances[10].u_tree.pipeline_current_node[0][7] ),
    .C1(_1997_),
    .X(_1998_));
 sky130_fd_sc_hd__inv_2 _4641_ (.A(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .Y(_1999_));
 sky130_fd_sc_hd__o22a_2 _4642_ (.A1(_1165_),
    .A2(_1999_),
    .B1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B2(_1595_),
    .X(_2000_));
 sky130_fd_sc_hd__o21ai_2 _4643_ (.A1(_1579_),
    .A2(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .B1(_2000_),
    .Y(_2001_));
 sky130_fd_sc_hd__a22o_2 _4644_ (.A1(_1578_),
    .A2(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .B1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .B2(_1596_),
    .X(_2002_));
 sky130_fd_sc_hd__xnor2_2 _4645_ (.A(_1159_),
    .B(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .Y(_2003_));
 sky130_fd_sc_hd__nand2_2 _4646_ (.A(_1599_),
    .B(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .Y(_2004_));
 sky130_fd_sc_hd__or4bb_2 _4647_ (.A(_1994_),
    .B(_2002_),
    .C_N(_2003_),
    .D_N(_2004_),
    .X(_2005_));
 sky130_fd_sc_hd__a2bb2o_2 _4648_ (.A1_N(_1598_),
    .A2_N(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .B1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .B2(_1581_),
    .X(_2006_));
 sky130_fd_sc_hd__a221o_2 _4649_ (.A1(_1165_),
    .A2(_1999_),
    .B1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B2(_1595_),
    .C1(_2006_),
    .X(_2007_));
 sky130_fd_sc_hd__or4_2 _4650_ (.A(_1998_),
    .B(_2001_),
    .C(_2005_),
    .D(_2007_),
    .X(_2008_));
 sky130_fd_sc_hd__nand2_2 _4651_ (.A(\tree_instances[10].u_tree.read_enable ),
    .B(_2008_),
    .Y(_2009_));
 sky130_fd_sc_hd__buf_1 _4652_ (.A(_2009_),
    .X(_2010_));
 sky130_fd_sc_hd__nand2_2 _4653_ (.A(_1994_),
    .B(_2010_),
    .Y(_0194_));
 sky130_fd_sc_hd__or3_2 _4654_ (.A(\tree_instances[0].u_tree.tree_state[1] ),
    .B(\tree_instances[0].u_tree.tree_state[2] ),
    .C(_1818_),
    .X(_2011_));
 sky130_fd_sc_hd__buf_1 _4655_ (.A(_2011_),
    .X(_2012_));
 sky130_fd_sc_hd__and2_2 _4656_ (.A(_1627_),
    .B(_2012_),
    .X(_2013_));
 sky130_fd_sc_hd__buf_1 _4657_ (.A(_2013_),
    .X(_0195_));
 sky130_fd_sc_hd__and2_2 _4658_ (.A(_1637_),
    .B(_2012_),
    .X(_2014_));
 sky130_fd_sc_hd__buf_1 _4659_ (.A(_2014_),
    .X(_0196_));
 sky130_fd_sc_hd__and2_2 _4660_ (.A(_1638_),
    .B(_2012_),
    .X(_2015_));
 sky130_fd_sc_hd__buf_1 _4661_ (.A(_2015_),
    .X(_0197_));
 sky130_fd_sc_hd__and2_2 _4662_ (.A(_1633_),
    .B(_2012_),
    .X(_2016_));
 sky130_fd_sc_hd__buf_1 _4663_ (.A(_2016_),
    .X(_0198_));
 sky130_fd_sc_hd__and2_2 _4664_ (.A(_1639_),
    .B(_2012_),
    .X(_2017_));
 sky130_fd_sc_hd__buf_1 _4665_ (.A(_2017_),
    .X(_0199_));
 sky130_fd_sc_hd__and2_2 _4666_ (.A(_1623_),
    .B(_2012_),
    .X(_2018_));
 sky130_fd_sc_hd__buf_1 _4667_ (.A(_2018_),
    .X(_0200_));
 sky130_fd_sc_hd__and2_2 _4668_ (.A(_1636_),
    .B(_2012_),
    .X(_2019_));
 sky130_fd_sc_hd__buf_1 _4669_ (.A(_2019_),
    .X(_0201_));
 sky130_fd_sc_hd__and2_2 _4670_ (.A(_1634_),
    .B(_2011_),
    .X(_2020_));
 sky130_fd_sc_hd__buf_1 _4671_ (.A(_2020_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_2 _4672_ (.A0(\tree_instances[10].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1827_),
    .S(_0006_),
    .X(_2021_));
 sky130_fd_sc_hd__buf_1 _4673_ (.A(_2021_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_2 _4674_ (.A0(\tree_instances[10].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1830_),
    .S(_0006_),
    .X(_2022_));
 sky130_fd_sc_hd__buf_1 _4675_ (.A(_2022_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_2 _4676_ (.A0(\tree_instances[10].u_tree.pipeline_frame_id[0][2] ),
    .A1(_1832_),
    .S(_0006_),
    .X(_2023_));
 sky130_fd_sc_hd__buf_1 _4677_ (.A(_2023_),
    .X(_0205_));
 sky130_fd_sc_hd__mux2_2 _4678_ (.A0(\tree_instances[10].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1835_),
    .S(_0006_),
    .X(_2024_));
 sky130_fd_sc_hd__buf_1 _4679_ (.A(_2024_),
    .X(_0206_));
 sky130_fd_sc_hd__mux2_2 _4680_ (.A0(\tree_instances[10].u_tree.pipeline_frame_id[0][4] ),
    .A1(_1837_),
    .S(_0006_),
    .X(_2025_));
 sky130_fd_sc_hd__buf_1 _4681_ (.A(_2025_),
    .X(_0207_));
 sky130_fd_sc_hd__inv_2 _4682_ (.A(\tree_instances[10].u_tree.read_enable ),
    .Y(_2026_));
 sky130_fd_sc_hd__buf_1 _4683_ (.A(_2026_),
    .X(_2027_));
 sky130_fd_sc_hd__o21ba_2 _4684_ (.A1(\tree_instances[10].u_tree.tree_state[0] ),
    .A2(_1172_),
    .B1_N(\tree_instances[10].u_tree.tree_state[1] ),
    .X(_2028_));
 sky130_fd_sc_hd__or3_2 _4685_ (.A(\tree_instances[10].u_tree.tree_state[1] ),
    .B(\tree_instances[10].u_tree.tree_state[2] ),
    .C(_1819_),
    .X(_2029_));
 sky130_fd_sc_hd__buf_1 _4686_ (.A(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__o21ai_2 _4687_ (.A1(_2027_),
    .A2(_2028_),
    .B1(_2030_),
    .Y(_0208_));
 sky130_fd_sc_hd__mux2_2 _4688_ (.A0(\tree_instances[10].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[10].u_tree.pipeline_frame_id[0][0] ),
    .S(_1136_),
    .X(_2031_));
 sky130_fd_sc_hd__buf_1 _4689_ (.A(_2031_),
    .X(_0209_));
 sky130_fd_sc_hd__mux2_2 _4690_ (.A0(\tree_instances[10].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[10].u_tree.pipeline_frame_id[0][1] ),
    .S(_1136_),
    .X(_2032_));
 sky130_fd_sc_hd__buf_1 _4691_ (.A(_2032_),
    .X(_0210_));
 sky130_fd_sc_hd__mux2_2 _4692_ (.A0(\tree_instances[10].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[10].u_tree.pipeline_frame_id[0][2] ),
    .S(_1136_),
    .X(_2033_));
 sky130_fd_sc_hd__buf_1 _4693_ (.A(_2033_),
    .X(_0211_));
 sky130_fd_sc_hd__mux2_2 _4694_ (.A0(\tree_instances[10].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[10].u_tree.pipeline_frame_id[0][3] ),
    .S(_1136_),
    .X(_2034_));
 sky130_fd_sc_hd__buf_1 _4695_ (.A(_2034_),
    .X(_0212_));
 sky130_fd_sc_hd__mux2_2 _4696_ (.A0(\tree_instances[10].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[10].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[10].u_tree.tree_state[3] ),
    .X(_2035_));
 sky130_fd_sc_hd__buf_1 _4697_ (.A(_2035_),
    .X(_0213_));
 sky130_fd_sc_hd__mux2_2 _4698_ (.A0(\tree_instances[10].u_tree.prediction_out ),
    .A1(\tree_instances[10].u_tree.pipeline_prediction[0][0] ),
    .S(\tree_instances[10].u_tree.tree_state[3] ),
    .X(_2036_));
 sky130_fd_sc_hd__buf_1 _4699_ (.A(_2036_),
    .X(_0214_));
 sky130_fd_sc_hd__a22o_2 _4700_ (.A1(_1136_),
    .A2(_1991_),
    .B1(_1819_),
    .B2(\tree_instances[10].u_tree.ready_for_next ),
    .X(_0215_));
 sky130_fd_sc_hd__o2bb2a_2 _4701_ (.A1_N(_0829_),
    .A2_N(_0830_),
    .B1(_0010_),
    .B2(\tree_instances[12].u_tree.pipeline_valid[0] ),
    .X(_0216_));
 sky130_fd_sc_hd__nand2_2 _4702_ (.A(_1591_),
    .B(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .Y(_2037_));
 sky130_fd_sc_hd__or2_2 _4703_ (.A(_1590_),
    .B(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .X(_2038_));
 sky130_fd_sc_hd__nand2_2 _4704_ (.A(_1573_),
    .B(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .Y(_2039_));
 sky130_fd_sc_hd__or2_2 _4705_ (.A(\tree_instances[10].u_tree.pipeline_current_node[0][6] ),
    .B(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .X(_2040_));
 sky130_fd_sc_hd__a221o_2 _4706_ (.A1(_2037_),
    .A2(_2038_),
    .B1(_2039_),
    .B2(_2040_),
    .C1(_1997_),
    .X(_2041_));
 sky130_fd_sc_hd__o221a_2 _4707_ (.A1(_1609_),
    .A2(_1999_),
    .B1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .B2(_1596_),
    .C1(_2004_),
    .X(_2042_));
 sky130_fd_sc_hd__o22a_2 _4708_ (.A1(_1581_),
    .A2(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .B1(_1996_),
    .B2(_1157_),
    .X(_2043_));
 sky130_fd_sc_hd__o221a_2 _4709_ (.A1(_1606_),
    .A2(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .B1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .B2(_1586_),
    .C1(_2043_),
    .X(_2044_));
 sky130_fd_sc_hd__o2111a_2 _4710_ (.A1(_1607_),
    .A2(_1995_),
    .B1(\tree_instances[10].u_tree.u_tree_weight_rom.cache_valid ),
    .C1(_2044_),
    .D1(_2003_),
    .X(_2045_));
 sky130_fd_sc_hd__and4bb_2 _4711_ (.A_N(_2026_),
    .B_N(_2041_),
    .C(_2042_),
    .D(_2045_),
    .X(_2046_));
 sky130_fd_sc_hd__buf_1 _4712_ (.A(_2046_),
    .X(_2047_));
 sky130_fd_sc_hd__buf_1 _4713_ (.A(_2047_),
    .X(_2048_));
 sky130_fd_sc_hd__and2_2 _4714_ (.A(\tree_instances[10].u_tree.read_enable ),
    .B(_2008_),
    .X(_2049_));
 sky130_fd_sc_hd__buf_1 _4715_ (.A(_2049_),
    .X(_2050_));
 sky130_fd_sc_hd__buf_1 _4716_ (.A(_2050_),
    .X(_2051_));
 sky130_fd_sc_hd__a22o_2 _4717_ (.A1(_2027_),
    .A2(\tree_instances[10].u_tree.node_data[12] ),
    .B1(_2051_),
    .B2(\tree_instances[10].u_tree.u_tree_weight_rom.gen_tree_10.u_tree_rom.node_data[12] ),
    .X(_2052_));
 sky130_fd_sc_hd__a21o_2 _4718_ (.A1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_data[12] ),
    .A2(_2048_),
    .B1(_2052_),
    .X(_0217_));
 sky130_fd_sc_hd__buf_1 _4719_ (.A(_2049_),
    .X(_2053_));
 sky130_fd_sc_hd__buf_1 _4720_ (.A(_2053_),
    .X(_2054_));
 sky130_fd_sc_hd__mux2_2 _4721_ (.A0(_1591_),
    .A1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .S(_2010_),
    .X(_2055_));
 sky130_fd_sc_hd__buf_1 _4722_ (.A(_2055_),
    .X(_0219_));
 sky130_fd_sc_hd__mux2_2 _4723_ (.A0(_1607_),
    .A1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .S(_2010_),
    .X(_2056_));
 sky130_fd_sc_hd__buf_1 _4724_ (.A(_2056_),
    .X(_0220_));
 sky130_fd_sc_hd__mux2_2 _4725_ (.A0(_1613_),
    .A1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .S(_2010_),
    .X(_2057_));
 sky130_fd_sc_hd__buf_1 _4726_ (.A(_2057_),
    .X(_0221_));
 sky130_fd_sc_hd__mux2_2 _4727_ (.A0(_1615_),
    .A1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .S(_2010_),
    .X(_2058_));
 sky130_fd_sc_hd__buf_1 _4728_ (.A(_2058_),
    .X(_0222_));
 sky130_fd_sc_hd__mux2_2 _4729_ (.A0(_1608_),
    .A1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .S(_2010_),
    .X(_2059_));
 sky130_fd_sc_hd__buf_1 _4730_ (.A(_2059_),
    .X(_0223_));
 sky130_fd_sc_hd__mux2_2 _4731_ (.A0(_1614_),
    .A1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .S(_2010_),
    .X(_2060_));
 sky130_fd_sc_hd__buf_1 _4732_ (.A(_2060_),
    .X(_0224_));
 sky130_fd_sc_hd__mux2_2 _4733_ (.A0(_1610_),
    .A1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .S(_2010_),
    .X(_2061_));
 sky130_fd_sc_hd__buf_1 _4734_ (.A(_2061_),
    .X(_0225_));
 sky130_fd_sc_hd__mux2_2 _4735_ (.A0(_1604_),
    .A1(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .S(_2009_),
    .X(_2062_));
 sky130_fd_sc_hd__buf_1 _4736_ (.A(_2062_),
    .X(_0226_));
 sky130_fd_sc_hd__mux2_2 _4737_ (.A0(\tree_instances[10].u_tree.u_tree_weight_rom.cached_data[12] ),
    .A1(\tree_instances[10].u_tree.u_tree_weight_rom.gen_tree_10.u_tree_rom.node_data[12] ),
    .S(_2054_),
    .X(_2063_));
 sky130_fd_sc_hd__buf_1 _4738_ (.A(_2063_),
    .X(_0227_));
 sky130_fd_sc_hd__mux2_2 _4739_ (.A0(\tree_instances[11].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1827_),
    .S(_0008_),
    .X(_2064_));
 sky130_fd_sc_hd__buf_1 _4740_ (.A(_2064_),
    .X(_0228_));
 sky130_fd_sc_hd__mux2_2 _4741_ (.A0(\tree_instances[11].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1830_),
    .S(_0008_),
    .X(_2065_));
 sky130_fd_sc_hd__buf_1 _4742_ (.A(_2065_),
    .X(_0229_));
 sky130_fd_sc_hd__mux2_2 _4743_ (.A0(\tree_instances[11].u_tree.pipeline_frame_id[0][2] ),
    .A1(_1832_),
    .S(_0008_),
    .X(_2066_));
 sky130_fd_sc_hd__buf_1 _4744_ (.A(_2066_),
    .X(_0230_));
 sky130_fd_sc_hd__mux2_2 _4745_ (.A0(\tree_instances[11].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1835_),
    .S(_0008_),
    .X(_2067_));
 sky130_fd_sc_hd__buf_1 _4746_ (.A(_2067_),
    .X(_0231_));
 sky130_fd_sc_hd__mux2_2 _4747_ (.A0(\tree_instances[11].u_tree.pipeline_frame_id[0][4] ),
    .A1(_1837_),
    .S(_0008_),
    .X(_2068_));
 sky130_fd_sc_hd__buf_1 _4748_ (.A(_2068_),
    .X(_0232_));
 sky130_fd_sc_hd__mux2_2 _4749_ (.A0(\tree_instances[10].u_tree.current_node_data[12] ),
    .A1(\tree_instances[10].u_tree.node_data[12] ),
    .S(_1172_),
    .X(_2069_));
 sky130_fd_sc_hd__buf_1 _4750_ (.A(_2069_),
    .X(_0233_));
 sky130_fd_sc_hd__or3_2 _4751_ (.A(\tree_instances[11].u_tree.tree_state[2] ),
    .B(\tree_instances[11].u_tree.tree_state[1] ),
    .C(_1816_),
    .X(_2070_));
 sky130_fd_sc_hd__buf_1 _4752_ (.A(_2070_),
    .X(_2071_));
 sky130_fd_sc_hd__mux2_2 _4753_ (.A0(\tree_instances[11].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[11].u_tree.pipeline_frame_id[0][0] ),
    .S(\tree_instances[11].u_tree.tree_state[3] ),
    .X(_2072_));
 sky130_fd_sc_hd__buf_1 _4754_ (.A(_2072_),
    .X(_0234_));
 sky130_fd_sc_hd__mux2_2 _4755_ (.A0(\tree_instances[11].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[11].u_tree.pipeline_frame_id[0][1] ),
    .S(\tree_instances[11].u_tree.tree_state[3] ),
    .X(_2073_));
 sky130_fd_sc_hd__buf_1 _4756_ (.A(_2073_),
    .X(_0235_));
 sky130_fd_sc_hd__mux2_2 _4757_ (.A0(\tree_instances[11].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[11].u_tree.pipeline_frame_id[0][2] ),
    .S(\tree_instances[11].u_tree.tree_state[3] ),
    .X(_2074_));
 sky130_fd_sc_hd__buf_1 _4758_ (.A(_2074_),
    .X(_0236_));
 sky130_fd_sc_hd__mux2_2 _4759_ (.A0(\tree_instances[11].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[11].u_tree.pipeline_frame_id[0][3] ),
    .S(\tree_instances[11].u_tree.tree_state[3] ),
    .X(_2075_));
 sky130_fd_sc_hd__buf_1 _4760_ (.A(_2075_),
    .X(_0237_));
 sky130_fd_sc_hd__mux2_2 _4761_ (.A0(\tree_instances[11].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[11].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[11].u_tree.tree_state[3] ),
    .X(_2076_));
 sky130_fd_sc_hd__buf_1 _4762_ (.A(_2076_),
    .X(_0238_));
 sky130_fd_sc_hd__and2_2 _4763_ (.A(_1591_),
    .B(_2030_),
    .X(_2077_));
 sky130_fd_sc_hd__buf_1 _4764_ (.A(_2077_),
    .X(_0239_));
 sky130_fd_sc_hd__and2_2 _4765_ (.A(_1607_),
    .B(_2030_),
    .X(_2078_));
 sky130_fd_sc_hd__buf_1 _4766_ (.A(_2078_),
    .X(_0240_));
 sky130_fd_sc_hd__and2_2 _4767_ (.A(_1613_),
    .B(_2030_),
    .X(_2079_));
 sky130_fd_sc_hd__buf_1 _4768_ (.A(_2079_),
    .X(_0241_));
 sky130_fd_sc_hd__and2_2 _4769_ (.A(_1615_),
    .B(_2030_),
    .X(_2080_));
 sky130_fd_sc_hd__buf_1 _4770_ (.A(_2080_),
    .X(_0242_));
 sky130_fd_sc_hd__and2_2 _4771_ (.A(_1608_),
    .B(_2030_),
    .X(_2081_));
 sky130_fd_sc_hd__buf_1 _4772_ (.A(_2081_),
    .X(_0243_));
 sky130_fd_sc_hd__and2_2 _4773_ (.A(_1614_),
    .B(_2030_),
    .X(_2082_));
 sky130_fd_sc_hd__buf_1 _4774_ (.A(_2082_),
    .X(_0244_));
 sky130_fd_sc_hd__and2_2 _4775_ (.A(_1610_),
    .B(_2030_),
    .X(_2083_));
 sky130_fd_sc_hd__buf_1 _4776_ (.A(_2083_),
    .X(_0245_));
 sky130_fd_sc_hd__and2_2 _4777_ (.A(_1604_),
    .B(_2029_),
    .X(_2084_));
 sky130_fd_sc_hd__buf_1 _4778_ (.A(_2084_),
    .X(_0246_));
 sky130_fd_sc_hd__a22o_2 _4779_ (.A1(\tree_instances[11].u_tree.tree_state[3] ),
    .A2(_0952_),
    .B1(_1816_),
    .B2(\tree_instances[11].u_tree.ready_for_next ),
    .X(_0247_));
 sky130_fd_sc_hd__and2_2 _4780_ (.A(_1429_),
    .B(_1430_),
    .X(_2085_));
 sky130_fd_sc_hd__buf_1 _4781_ (.A(_2085_),
    .X(_0248_));
 sky130_fd_sc_hd__buf_1 _4782_ (.A(\tree_instances[12].u_tree.tree_state[2] ),
    .X(_2086_));
 sky130_fd_sc_hd__a22o_2 _4783_ (.A1(\tree_instances[12].u_tree.tree_state[1] ),
    .A2(\tree_instances[12].u_tree.current_node_data[12] ),
    .B1(\tree_instances[12].u_tree.node_data[12] ),
    .B2(_2086_),
    .X(_2087_));
 sky130_fd_sc_hd__o31ai_2 _4784_ (.A1(\tree_instances[12].u_tree.tree_state[0] ),
    .A2(\tree_instances[12].u_tree.tree_state[1] ),
    .A3(\tree_instances[12].u_tree.tree_state[2] ),
    .B1(_0830_),
    .Y(_2088_));
 sky130_fd_sc_hd__or2_2 _4785_ (.A(_0009_),
    .B(_2088_),
    .X(_2089_));
 sky130_fd_sc_hd__mux2_2 _4786_ (.A0(_2087_),
    .A1(\tree_instances[12].u_tree.pipeline_prediction[0][0] ),
    .S(_2089_),
    .X(_2090_));
 sky130_fd_sc_hd__buf_1 _4787_ (.A(_2090_),
    .X(_0249_));
 sky130_fd_sc_hd__inv_2 _4788_ (.A(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .Y(_2091_));
 sky130_fd_sc_hd__a22o_2 _4789_ (.A1(_1702_),
    .A2(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .B1(_2091_),
    .B2(_0839_),
    .X(_2092_));
 sky130_fd_sc_hd__a221o_2 _4790_ (.A1(_1711_),
    .A2(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .B1(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .B2(_1691_),
    .C1(_2092_),
    .X(_2093_));
 sky130_fd_sc_hd__or2_2 _4791_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][7] ),
    .B(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .X(_2094_));
 sky130_fd_sc_hd__nand2_2 _4792_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][7] ),
    .B(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .Y(_2095_));
 sky130_fd_sc_hd__nand2_2 _4793_ (.A(_0838_),
    .B(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .Y(_2096_));
 sky130_fd_sc_hd__or2_2 _4794_ (.A(_0837_),
    .B(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .X(_2097_));
 sky130_fd_sc_hd__xor2_2 _4795_ (.A(\tree_instances[12].u_tree.pipeline_current_node[0][6] ),
    .B(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .X(_2098_));
 sky130_fd_sc_hd__a221o_2 _4796_ (.A1(_2094_),
    .A2(_2095_),
    .B1(_2096_),
    .B2(_2097_),
    .C1(_2098_),
    .X(_2099_));
 sky130_fd_sc_hd__or2_2 _4797_ (.A(_1698_),
    .B(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .X(_2100_));
 sky130_fd_sc_hd__or2_2 _4798_ (.A(_1711_),
    .B(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .X(_2101_));
 sky130_fd_sc_hd__or2_2 _4799_ (.A(_0839_),
    .B(_2091_),
    .X(_2102_));
 sky130_fd_sc_hd__and3_2 _4800_ (.A(_2100_),
    .B(_2101_),
    .C(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__or2_2 _4801_ (.A(_1691_),
    .B(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .X(_2104_));
 sky130_fd_sc_hd__or2_2 _4802_ (.A(_1702_),
    .B(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .X(_2105_));
 sky130_fd_sc_hd__nand2_2 _4803_ (.A(_1698_),
    .B(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .Y(_2106_));
 sky130_fd_sc_hd__and4_2 _4804_ (.A(\tree_instances[12].u_tree.u_tree_weight_rom.cache_valid ),
    .B(_2104_),
    .C(_2105_),
    .D(_2106_),
    .X(_2107_));
 sky130_fd_sc_hd__or4bb_2 _4805_ (.A(_2093_),
    .B(_2099_),
    .C_N(_2103_),
    .D_N(_2107_),
    .X(_2108_));
 sky130_fd_sc_hd__and2_2 _4806_ (.A(\tree_instances[12].u_tree.read_enable ),
    .B(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__buf_1 _4807_ (.A(_2109_),
    .X(_2110_));
 sky130_fd_sc_hd__buf_1 _4808_ (.A(_2110_),
    .X(_2111_));
 sky130_fd_sc_hd__buf_1 _4809_ (.A(_2111_),
    .X(_2112_));
 sky130_fd_sc_hd__or2_2 _4810_ (.A(\tree_instances[12].u_tree.u_tree_weight_rom.cache_valid ),
    .B(_2112_),
    .X(_2113_));
 sky130_fd_sc_hd__buf_1 _4811_ (.A(_2113_),
    .X(_0250_));
 sky130_fd_sc_hd__and2_2 _4812_ (.A(_1275_),
    .B(_2071_),
    .X(_2114_));
 sky130_fd_sc_hd__buf_1 _4813_ (.A(_2114_),
    .X(_0251_));
 sky130_fd_sc_hd__and2_2 _4814_ (.A(_1276_),
    .B(_2071_),
    .X(_2115_));
 sky130_fd_sc_hd__buf_1 _4815_ (.A(_2115_),
    .X(_0252_));
 sky130_fd_sc_hd__and2_2 _4816_ (.A(_1274_),
    .B(_2071_),
    .X(_2116_));
 sky130_fd_sc_hd__buf_1 _4817_ (.A(_2116_),
    .X(_0253_));
 sky130_fd_sc_hd__and2_2 _4818_ (.A(_1278_),
    .B(_2071_),
    .X(_2117_));
 sky130_fd_sc_hd__buf_1 _4819_ (.A(_2117_),
    .X(_0254_));
 sky130_fd_sc_hd__and2_2 _4820_ (.A(_1284_),
    .B(_2071_),
    .X(_2118_));
 sky130_fd_sc_hd__buf_1 _4821_ (.A(_2118_),
    .X(_0255_));
 sky130_fd_sc_hd__and2_2 _4822_ (.A(_1281_),
    .B(_2071_),
    .X(_2119_));
 sky130_fd_sc_hd__buf_1 _4823_ (.A(_2119_),
    .X(_0256_));
 sky130_fd_sc_hd__and2_2 _4824_ (.A(_1286_),
    .B(_2071_),
    .X(_2120_));
 sky130_fd_sc_hd__buf_1 _4825_ (.A(_2120_),
    .X(_0257_));
 sky130_fd_sc_hd__and2_2 _4826_ (.A(_1285_),
    .B(_2070_),
    .X(_2121_));
 sky130_fd_sc_hd__buf_1 _4827_ (.A(_2121_),
    .X(_0258_));
 sky130_fd_sc_hd__buf_1 _4828_ (.A(\tree_instances[0].u_tree.frame_id_in[0] ),
    .X(_2122_));
 sky130_fd_sc_hd__mux2_2 _4829_ (.A0(\tree_instances[12].u_tree.pipeline_frame_id[0][0] ),
    .A1(_2122_),
    .S(_0010_),
    .X(_2123_));
 sky130_fd_sc_hd__buf_1 _4830_ (.A(_2123_),
    .X(_0259_));
 sky130_fd_sc_hd__mux2_2 _4831_ (.A0(\tree_instances[12].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1830_),
    .S(_0010_),
    .X(_2124_));
 sky130_fd_sc_hd__buf_1 _4832_ (.A(_2124_),
    .X(_0260_));
 sky130_fd_sc_hd__buf_1 _4833_ (.A(\tree_instances[0].u_tree.frame_id_in[2] ),
    .X(_2125_));
 sky130_fd_sc_hd__mux2_2 _4834_ (.A0(\tree_instances[12].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2125_),
    .S(_0010_),
    .X(_2126_));
 sky130_fd_sc_hd__buf_1 _4835_ (.A(_2126_),
    .X(_0261_));
 sky130_fd_sc_hd__mux2_2 _4836_ (.A0(\tree_instances[12].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1835_),
    .S(_0010_),
    .X(_2127_));
 sky130_fd_sc_hd__buf_1 _4837_ (.A(_2127_),
    .X(_0262_));
 sky130_fd_sc_hd__mux2_2 _4838_ (.A0(\tree_instances[12].u_tree.pipeline_frame_id[0][4] ),
    .A1(_1837_),
    .S(_0010_),
    .X(_2128_));
 sky130_fd_sc_hd__buf_1 _4839_ (.A(_2128_),
    .X(_0263_));
 sky130_fd_sc_hd__inv_2 _4840_ (.A(\tree_instances[12].u_tree.read_enable ),
    .Y(_2129_));
 sky130_fd_sc_hd__buf_1 _4841_ (.A(_2129_),
    .X(_2130_));
 sky130_fd_sc_hd__o21ba_2 _4842_ (.A1(\tree_instances[12].u_tree.tree_state[0] ),
    .A2(_1026_),
    .B1_N(\tree_instances[12].u_tree.tree_state[1] ),
    .X(_2131_));
 sky130_fd_sc_hd__or3_2 _4843_ (.A(\tree_instances[12].u_tree.tree_state[1] ),
    .B(\tree_instances[12].u_tree.tree_state[2] ),
    .C(_1810_),
    .X(_2132_));
 sky130_fd_sc_hd__buf_1 _4844_ (.A(_2132_),
    .X(_2133_));
 sky130_fd_sc_hd__o21ai_2 _4845_ (.A1(_2130_),
    .A2(_2131_),
    .B1(_2133_),
    .Y(_0264_));
 sky130_fd_sc_hd__mux2_2 _4846_ (.A0(\tree_instances[12].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[12].u_tree.pipeline_frame_id[0][0] ),
    .S(_0829_),
    .X(_2134_));
 sky130_fd_sc_hd__buf_1 _4847_ (.A(_2134_),
    .X(_0265_));
 sky130_fd_sc_hd__mux2_2 _4848_ (.A0(\tree_instances[12].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[12].u_tree.pipeline_frame_id[0][1] ),
    .S(_0829_),
    .X(_2135_));
 sky130_fd_sc_hd__buf_1 _4849_ (.A(_2135_),
    .X(_0266_));
 sky130_fd_sc_hd__mux2_2 _4850_ (.A0(\tree_instances[12].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[12].u_tree.pipeline_frame_id[0][2] ),
    .S(_0829_),
    .X(_2136_));
 sky130_fd_sc_hd__buf_1 _4851_ (.A(_2136_),
    .X(_0267_));
 sky130_fd_sc_hd__mux2_2 _4852_ (.A0(\tree_instances[12].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[12].u_tree.pipeline_frame_id[0][3] ),
    .S(_0829_),
    .X(_2137_));
 sky130_fd_sc_hd__buf_1 _4853_ (.A(_2137_),
    .X(_0268_));
 sky130_fd_sc_hd__mux2_2 _4854_ (.A0(\tree_instances[12].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[12].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[12].u_tree.tree_state[3] ),
    .X(_2138_));
 sky130_fd_sc_hd__buf_1 _4855_ (.A(_2138_),
    .X(_0269_));
 sky130_fd_sc_hd__mux2_2 _4856_ (.A0(\tree_instances[12].u_tree.prediction_out ),
    .A1(\tree_instances[12].u_tree.pipeline_prediction[0][0] ),
    .S(\tree_instances[12].u_tree.tree_state[3] ),
    .X(_2139_));
 sky130_fd_sc_hd__buf_1 _4857_ (.A(_2139_),
    .X(_0270_));
 sky130_fd_sc_hd__a22o_2 _4858_ (.A1(_0829_),
    .A2(_0830_),
    .B1(_1810_),
    .B2(\tree_instances[12].u_tree.ready_for_next ),
    .X(_0271_));
 sky130_fd_sc_hd__buf_1 _4859_ (.A(_0825_),
    .X(_2140_));
 sky130_fd_sc_hd__buf_1 _4860_ (.A(_0823_),
    .X(_2141_));
 sky130_fd_sc_hd__buf_1 _4861_ (.A(_2141_),
    .X(_2142_));
 sky130_fd_sc_hd__buf_1 _4862_ (.A(_0821_),
    .X(_2143_));
 sky130_fd_sc_hd__buf_1 _4863_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][1] ),
    .X(_2144_));
 sky130_fd_sc_hd__buf_1 _4864_ (.A(_2144_),
    .X(_2145_));
 sky130_fd_sc_hd__buf_1 _4865_ (.A(_0813_),
    .X(_2146_));
 sky130_fd_sc_hd__buf_1 _4866_ (.A(_2142_),
    .X(_2147_));
 sky130_fd_sc_hd__buf_1 _4867_ (.A(_2143_),
    .X(_2148_));
 sky130_fd_sc_hd__buf_1 _4868_ (.A(_2145_),
    .X(_2149_));
 sky130_fd_sc_hd__buf_1 _4869_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][7] ),
    .X(_2150_));
 sky130_fd_sc_hd__buf_1 _4870_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][8] ),
    .X(_2151_));
 sky130_fd_sc_hd__buf_1 _4871_ (.A(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__buf_1 _4872_ (.A(_0810_),
    .X(_2153_));
 sky130_fd_sc_hd__buf_1 _4873_ (.A(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__buf_1 _4874_ (.A(_2146_),
    .X(_2155_));
 sky130_fd_sc_hd__buf_1 _4875_ (.A(_0818_),
    .X(_2156_));
 sky130_fd_sc_hd__buf_1 _4876_ (.A(_2156_),
    .X(_2157_));
 sky130_fd_sc_hd__buf_1 _4877_ (.A(_2140_),
    .X(_2158_));
 sky130_fd_sc_hd__buf_1 _4878_ (.A(_2150_),
    .X(_2159_));
 sky130_fd_sc_hd__buf_1 _4879_ (.A(_2154_),
    .X(_2160_));
 sky130_fd_sc_hd__buf_1 _4880_ (.A(_2148_),
    .X(_2161_));
 sky130_fd_sc_hd__buf_1 _4881_ (.A(_2155_),
    .X(_2162_));
 sky130_fd_sc_hd__buf_1 _4882_ (.A(_2158_),
    .X(_2163_));
 sky130_fd_sc_hd__buf_1 _4883_ (.A(_0967_),
    .X(_2164_));
 sky130_fd_sc_hd__a22o_2 _4884_ (.A1(\tree_instances[13].u_tree.tree_state[1] ),
    .A2(\tree_instances[13].u_tree.current_node_data[12] ),
    .B1(\tree_instances[13].u_tree.node_data[12] ),
    .B2(_2164_),
    .X(_2165_));
 sky130_fd_sc_hd__nor3_2 _4885_ (.A(\tree_instances[13].u_tree.tree_state[1] ),
    .B(_0967_),
    .C(\tree_instances[13].u_tree.tree_state[0] ),
    .Y(_2166_));
 sky130_fd_sc_hd__a211o_2 _4886_ (.A1(\tree_instances[13].u_tree.tree_state[0] ),
    .A2(_1113_),
    .B1(_2166_),
    .C1(_0011_),
    .X(_2167_));
 sky130_fd_sc_hd__mux2_2 _4887_ (.A0(_2165_),
    .A1(\tree_instances[13].u_tree.pipeline_prediction[0][0] ),
    .S(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__buf_1 _4888_ (.A(_2168_),
    .X(_0272_));
 sky130_fd_sc_hd__inv_2 _4889_ (.A(\tree_instances[13].u_tree.u_tree_weight_rom.cache_valid ),
    .Y(_2169_));
 sky130_fd_sc_hd__inv_2 _4890_ (.A(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .Y(_2170_));
 sky130_fd_sc_hd__xor2_2 _4891_ (.A(_1650_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .X(_2171_));
 sky130_fd_sc_hd__nand2_2 _4892_ (.A(_0953_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .Y(_2172_));
 sky130_fd_sc_hd__or2_2 _4893_ (.A(_0953_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .X(_2173_));
 sky130_fd_sc_hd__nand2_2 _4894_ (.A(_2172_),
    .B(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__nor2_2 _4895_ (.A(_1656_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .Y(_2175_));
 sky130_fd_sc_hd__and2_2 _4896_ (.A(_0962_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .X(_2176_));
 sky130_fd_sc_hd__a2111o_2 _4897_ (.A1(_1654_),
    .A2(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .B1(_2169_),
    .C1(_2175_),
    .D1(_2176_),
    .X(_2177_));
 sky130_fd_sc_hd__and2_2 _4898_ (.A(_1640_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .X(_2178_));
 sky130_fd_sc_hd__nor2_2 _4899_ (.A(_0963_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .Y(_2179_));
 sky130_fd_sc_hd__o21bai_2 _4900_ (.A1(_1662_),
    .A2(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B1_N(_2179_),
    .Y(_2180_));
 sky130_fd_sc_hd__a211o_2 _4901_ (.A1(_1662_),
    .A2(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B1(_2178_),
    .C1(_2180_),
    .X(_2181_));
 sky130_fd_sc_hd__and2_2 _4902_ (.A(_1656_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .X(_2182_));
 sky130_fd_sc_hd__and2b_2 _4903_ (.A_N(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .B(_0958_),
    .X(_2183_));
 sky130_fd_sc_hd__and2b_2 _4904_ (.A_N(_0958_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .X(_2184_));
 sky130_fd_sc_hd__nor2_2 _4905_ (.A(_1641_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .Y(_2185_));
 sky130_fd_sc_hd__or4_2 _4906_ (.A(_2182_),
    .B(_2183_),
    .C(_2184_),
    .D(_2185_),
    .X(_2186_));
 sky130_fd_sc_hd__or4_2 _4907_ (.A(_2174_),
    .B(_2177_),
    .C(_2181_),
    .D(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__a211o_2 _4908_ (.A1(_1686_),
    .A2(_2170_),
    .B1(_2171_),
    .C1(_2187_),
    .X(_2188_));
 sky130_fd_sc_hd__nand2_2 _4909_ (.A(\tree_instances[13].u_tree.read_enable ),
    .B(_2188_),
    .Y(_2189_));
 sky130_fd_sc_hd__buf_1 _4910_ (.A(_2189_),
    .X(_2190_));
 sky130_fd_sc_hd__buf_1 _4911_ (.A(_2190_),
    .X(_2191_));
 sky130_fd_sc_hd__nand2_2 _4912_ (.A(_2169_),
    .B(_2191_),
    .Y(_0273_));
 sky130_fd_sc_hd__nand2_2 _4913_ (.A(\tree_instances[12].u_tree.read_enable ),
    .B(_2108_),
    .Y(_2192_));
 sky130_fd_sc_hd__mux2_2 _4914_ (.A0(_1708_),
    .A1(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .S(_2192_),
    .X(_2193_));
 sky130_fd_sc_hd__buf_1 _4915_ (.A(_2193_),
    .X(_0274_));
 sky130_fd_sc_hd__mux2_2 _4916_ (.A0(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .A1(_1713_),
    .S(\tree_instances[12].u_tree.read_enable ),
    .X(_2194_));
 sky130_fd_sc_hd__buf_1 _4917_ (.A(_2194_),
    .X(_0275_));
 sky130_fd_sc_hd__mux2_2 _4918_ (.A0(_1723_),
    .A1(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .S(_2192_),
    .X(_2195_));
 sky130_fd_sc_hd__buf_1 _4919_ (.A(_2195_),
    .X(_0276_));
 sky130_fd_sc_hd__mux2_2 _4920_ (.A0(_1724_),
    .A1(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .S(_2192_),
    .X(_2196_));
 sky130_fd_sc_hd__buf_1 _4921_ (.A(_2196_),
    .X(_0277_));
 sky130_fd_sc_hd__mux2_2 _4922_ (.A0(_1727_),
    .A1(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .S(_2192_),
    .X(_2197_));
 sky130_fd_sc_hd__buf_1 _4923_ (.A(_2197_),
    .X(_0278_));
 sky130_fd_sc_hd__mux2_2 _4924_ (.A0(_1721_),
    .A1(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .S(_2192_),
    .X(_2198_));
 sky130_fd_sc_hd__buf_1 _4925_ (.A(_2198_),
    .X(_0279_));
 sky130_fd_sc_hd__mux2_2 _4926_ (.A0(_1726_),
    .A1(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .S(_2192_),
    .X(_2199_));
 sky130_fd_sc_hd__buf_1 _4927_ (.A(_2199_),
    .X(_0280_));
 sky130_fd_sc_hd__mux2_2 _4928_ (.A0(_1718_),
    .A1(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .S(_2192_),
    .X(_2200_));
 sky130_fd_sc_hd__buf_1 _4929_ (.A(_2200_),
    .X(_0281_));
 sky130_fd_sc_hd__buf_1 _4930_ (.A(_2111_),
    .X(_2201_));
 sky130_fd_sc_hd__mux2_2 _4931_ (.A0(\tree_instances[12].u_tree.u_tree_weight_rom.cached_data[12] ),
    .A1(\tree_instances[12].u_tree.u_tree_weight_rom.gen_tree_12.u_tree_rom.node_data[12] ),
    .S(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__buf_1 _4932_ (.A(_2202_),
    .X(_0282_));
 sky130_fd_sc_hd__and3_2 _4933_ (.A(_1673_),
    .B(_1683_),
    .C(_1685_),
    .X(_2203_));
 sky130_fd_sc_hd__buf_1 _4934_ (.A(_2203_),
    .X(_0283_));
 sky130_fd_sc_hd__and2_2 _4935_ (.A(_1708_),
    .B(_2133_),
    .X(_2204_));
 sky130_fd_sc_hd__buf_1 _4936_ (.A(_2204_),
    .X(_0284_));
 sky130_fd_sc_hd__and2_2 _4937_ (.A(_1713_),
    .B(_2133_),
    .X(_2205_));
 sky130_fd_sc_hd__buf_1 _4938_ (.A(_2205_),
    .X(_0285_));
 sky130_fd_sc_hd__and2_2 _4939_ (.A(_1723_),
    .B(_2133_),
    .X(_2206_));
 sky130_fd_sc_hd__buf_1 _4940_ (.A(_2206_),
    .X(_0286_));
 sky130_fd_sc_hd__and2_2 _4941_ (.A(_1724_),
    .B(_2133_),
    .X(_2207_));
 sky130_fd_sc_hd__buf_1 _4942_ (.A(_2207_),
    .X(_0287_));
 sky130_fd_sc_hd__and2_2 _4943_ (.A(_1727_),
    .B(_2133_),
    .X(_2208_));
 sky130_fd_sc_hd__buf_1 _4944_ (.A(_2208_),
    .X(_0288_));
 sky130_fd_sc_hd__and2_2 _4945_ (.A(_1721_),
    .B(_2133_),
    .X(_2209_));
 sky130_fd_sc_hd__buf_1 _4946_ (.A(_2209_),
    .X(_0289_));
 sky130_fd_sc_hd__and2_2 _4947_ (.A(_1726_),
    .B(_2133_),
    .X(_2210_));
 sky130_fd_sc_hd__buf_1 _4948_ (.A(_2210_),
    .X(_0290_));
 sky130_fd_sc_hd__and2_2 _4949_ (.A(_1718_),
    .B(_2132_),
    .X(_2211_));
 sky130_fd_sc_hd__buf_1 _4950_ (.A(_2211_),
    .X(_0291_));
 sky130_fd_sc_hd__mux2_2 _4951_ (.A0(_1827_),
    .A1(\tree_instances[13].u_tree.pipeline_frame_id[0][0] ),
    .S(_1824_),
    .X(_2212_));
 sky130_fd_sc_hd__buf_1 _4952_ (.A(_2212_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_2 _4953_ (.A0(_1830_),
    .A1(\tree_instances[13].u_tree.pipeline_frame_id[0][1] ),
    .S(_1824_),
    .X(_2213_));
 sky130_fd_sc_hd__buf_1 _4954_ (.A(_2213_),
    .X(_0293_));
 sky130_fd_sc_hd__mux2_2 _4955_ (.A0(_1832_),
    .A1(\tree_instances[13].u_tree.pipeline_frame_id[0][2] ),
    .S(_1824_),
    .X(_2214_));
 sky130_fd_sc_hd__buf_1 _4956_ (.A(_2214_),
    .X(_0294_));
 sky130_fd_sc_hd__mux2_2 _4957_ (.A0(_1835_),
    .A1(\tree_instances[13].u_tree.pipeline_frame_id[0][3] ),
    .S(_1824_),
    .X(_2215_));
 sky130_fd_sc_hd__buf_1 _4958_ (.A(_2215_),
    .X(_0295_));
 sky130_fd_sc_hd__mux2_2 _4959_ (.A0(_1837_),
    .A1(\tree_instances[13].u_tree.pipeline_frame_id[0][4] ),
    .S(_1824_),
    .X(_2216_));
 sky130_fd_sc_hd__buf_1 _4960_ (.A(_2216_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_2 _4961_ (.A0(\tree_instances[12].u_tree.current_node_data[12] ),
    .A1(\tree_instances[12].u_tree.node_data[12] ),
    .S(_1026_),
    .X(_2217_));
 sky130_fd_sc_hd__buf_1 _4962_ (.A(_2217_),
    .X(_0297_));
 sky130_fd_sc_hd__inv_2 _4963_ (.A(\tree_instances[13].u_tree.read_enable ),
    .Y(_2218_));
 sky130_fd_sc_hd__buf_1 _4964_ (.A(_2218_),
    .X(_2219_));
 sky130_fd_sc_hd__nor2_2 _4965_ (.A(\tree_instances[13].u_tree.tree_state[1] ),
    .B(_2166_),
    .Y(_2220_));
 sky130_fd_sc_hd__or3_2 _4966_ (.A(\tree_instances[13].u_tree.tree_state[1] ),
    .B(_0967_),
    .C(_1823_),
    .X(_2221_));
 sky130_fd_sc_hd__buf_1 _4967_ (.A(_2221_),
    .X(_2222_));
 sky130_fd_sc_hd__o21ai_2 _4968_ (.A1(_2219_),
    .A2(_2220_),
    .B1(_2222_),
    .Y(_0298_));
 sky130_fd_sc_hd__mux2_2 _4969_ (.A0(\tree_instances[13].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[13].u_tree.pipeline_frame_id[0][0] ),
    .S(_1114_),
    .X(_2223_));
 sky130_fd_sc_hd__buf_1 _4970_ (.A(_2223_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_2 _4971_ (.A0(\tree_instances[13].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[13].u_tree.pipeline_frame_id[0][1] ),
    .S(_1114_),
    .X(_2224_));
 sky130_fd_sc_hd__buf_1 _4972_ (.A(_2224_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_2 _4973_ (.A0(\tree_instances[13].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[13].u_tree.pipeline_frame_id[0][2] ),
    .S(_1114_),
    .X(_2225_));
 sky130_fd_sc_hd__buf_1 _4974_ (.A(_2225_),
    .X(_0301_));
 sky130_fd_sc_hd__mux2_2 _4975_ (.A0(\tree_instances[13].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[13].u_tree.pipeline_frame_id[0][3] ),
    .S(\tree_instances[13].u_tree.tree_state[3] ),
    .X(_2226_));
 sky130_fd_sc_hd__buf_1 _4976_ (.A(_2226_),
    .X(_0302_));
 sky130_fd_sc_hd__mux2_2 _4977_ (.A0(\tree_instances[13].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[13].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[13].u_tree.tree_state[3] ),
    .X(_2227_));
 sky130_fd_sc_hd__buf_1 _4978_ (.A(_2227_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_2 _4979_ (.A0(\tree_instances[13].u_tree.prediction_out ),
    .A1(\tree_instances[13].u_tree.pipeline_prediction[0][0] ),
    .S(\tree_instances[13].u_tree.tree_state[3] ),
    .X(_2228_));
 sky130_fd_sc_hd__buf_1 _4980_ (.A(_2228_),
    .X(_0304_));
 sky130_fd_sc_hd__a21oi_2 _4981_ (.A1(_1822_),
    .A2(_1114_),
    .B1(\tree_instances[13].u_tree.ready_for_next ),
    .Y(_2229_));
 sky130_fd_sc_hd__nor2_2 _4982_ (.A(_1114_),
    .B(_1824_),
    .Y(_2230_));
 sky130_fd_sc_hd__a21oi_2 _4983_ (.A1(_1824_),
    .A2(_2229_),
    .B1(_2230_),
    .Y(_0305_));
 sky130_fd_sc_hd__o2bb2a_2 _4984_ (.A1_N(_1822_),
    .A2_N(_1114_),
    .B1(_2230_),
    .B2(\tree_instances[13].u_tree.pipeline_valid[0] ),
    .X(_0306_));
 sky130_fd_sc_hd__buf_1 _4985_ (.A(_2189_),
    .X(_2231_));
 sky130_fd_sc_hd__mux2_2 _4986_ (.A0(_1666_),
    .A1(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .S(_2231_),
    .X(_2232_));
 sky130_fd_sc_hd__buf_1 _4987_ (.A(_2232_),
    .X(_0307_));
 sky130_fd_sc_hd__mux2_2 _4988_ (.A0(_1679_),
    .A1(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .S(_2231_),
    .X(_2233_));
 sky130_fd_sc_hd__buf_1 _4989_ (.A(_2233_),
    .X(_0308_));
 sky130_fd_sc_hd__mux2_2 _4990_ (.A0(_1686_),
    .A1(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .S(_2231_),
    .X(_2234_));
 sky130_fd_sc_hd__buf_1 _4991_ (.A(_2234_),
    .X(_0309_));
 sky130_fd_sc_hd__mux2_2 _4992_ (.A0(_1684_),
    .A1(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .S(_2231_),
    .X(_2235_));
 sky130_fd_sc_hd__buf_1 _4993_ (.A(_2235_),
    .X(_0310_));
 sky130_fd_sc_hd__mux2_2 _4994_ (.A0(_1647_),
    .A1(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .S(_2189_),
    .X(_2236_));
 sky130_fd_sc_hd__buf_1 _4995_ (.A(_2236_),
    .X(_0311_));
 sky130_fd_sc_hd__mux2_2 _4996_ (.A0(_1676_),
    .A1(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .S(_2189_),
    .X(_2237_));
 sky130_fd_sc_hd__buf_1 _4997_ (.A(_2237_),
    .X(_0312_));
 sky130_fd_sc_hd__mux2_2 _4998_ (.A0(_1669_),
    .A1(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .S(_2189_),
    .X(_2238_));
 sky130_fd_sc_hd__buf_1 _4999_ (.A(_2238_),
    .X(_0313_));
 sky130_fd_sc_hd__mux2_2 _5000_ (.A0(_1673_),
    .A1(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .S(_2189_),
    .X(_2239_));
 sky130_fd_sc_hd__buf_1 _5001_ (.A(_2239_),
    .X(_0314_));
 sky130_fd_sc_hd__buf_1 _5002_ (.A(\tree_instances[13].u_tree.read_enable ),
    .X(_2240_));
 sky130_fd_sc_hd__buf_1 _5003_ (.A(_2240_),
    .X(_2241_));
 sky130_fd_sc_hd__buf_1 _5004_ (.A(_2188_),
    .X(_2242_));
 sky130_fd_sc_hd__buf_1 _5005_ (.A(_2242_),
    .X(_2243_));
 sky130_fd_sc_hd__and3_2 _5006_ (.A(_2241_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.gen_tree_13.u_tree_rom.node_data[12] ),
    .C(_2243_),
    .X(_2244_));
 sky130_fd_sc_hd__a21o_2 _5007_ (.A1(\tree_instances[13].u_tree.u_tree_weight_rom.cached_data[12] ),
    .A2(_2191_),
    .B1(_2244_),
    .X(_0315_));
 sky130_fd_sc_hd__mux2_2 _5008_ (.A0(\tree_instances[14].u_tree.pipeline_frame_id[0][0] ),
    .A1(_2122_),
    .S(_0014_),
    .X(_2245_));
 sky130_fd_sc_hd__buf_1 _5009_ (.A(_2245_),
    .X(_0316_));
 sky130_fd_sc_hd__buf_1 _5010_ (.A(_1829_),
    .X(_2246_));
 sky130_fd_sc_hd__mux2_2 _5011_ (.A0(\tree_instances[14].u_tree.pipeline_frame_id[0][1] ),
    .A1(_2246_),
    .S(_0014_),
    .X(_2247_));
 sky130_fd_sc_hd__buf_1 _5012_ (.A(_2247_),
    .X(_0317_));
 sky130_fd_sc_hd__mux2_2 _5013_ (.A0(\tree_instances[14].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2125_),
    .S(_0014_),
    .X(_2248_));
 sky130_fd_sc_hd__buf_1 _5014_ (.A(_2248_),
    .X(_0318_));
 sky130_fd_sc_hd__buf_1 _5015_ (.A(\tree_instances[0].u_tree.frame_id_in[3] ),
    .X(_2249_));
 sky130_fd_sc_hd__mux2_2 _5016_ (.A0(\tree_instances[14].u_tree.pipeline_frame_id[0][3] ),
    .A1(_2249_),
    .S(_0014_),
    .X(_2250_));
 sky130_fd_sc_hd__buf_1 _5017_ (.A(_2250_),
    .X(_0319_));
 sky130_fd_sc_hd__buf_1 _5018_ (.A(\tree_instances[0].u_tree.frame_id_in[4] ),
    .X(_2251_));
 sky130_fd_sc_hd__mux2_2 _5019_ (.A0(\tree_instances[14].u_tree.pipeline_frame_id[0][4] ),
    .A1(_2251_),
    .S(_0014_),
    .X(_2252_));
 sky130_fd_sc_hd__buf_1 _5020_ (.A(_2252_),
    .X(_0320_));
 sky130_fd_sc_hd__mux2_2 _5021_ (.A0(\tree_instances[13].u_tree.current_node_data[12] ),
    .A1(\tree_instances[13].u_tree.node_data[12] ),
    .S(_0968_),
    .X(_2253_));
 sky130_fd_sc_hd__buf_1 _5022_ (.A(_2253_),
    .X(_0321_));
 sky130_fd_sc_hd__or3_2 _5023_ (.A(\tree_instances[14].u_tree.tree_state[1] ),
    .B(\tree_instances[14].u_tree.tree_state[2] ),
    .C(_1817_),
    .X(_2254_));
 sky130_fd_sc_hd__buf_1 _5024_ (.A(_2254_),
    .X(_2255_));
 sky130_fd_sc_hd__mux2_2 _5025_ (.A0(\tree_instances[14].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[14].u_tree.pipeline_frame_id[0][0] ),
    .S(_0735_),
    .X(_2256_));
 sky130_fd_sc_hd__buf_1 _5026_ (.A(_2256_),
    .X(_0322_));
 sky130_fd_sc_hd__mux2_2 _5027_ (.A0(\tree_instances[14].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[14].u_tree.pipeline_frame_id[0][1] ),
    .S(_0735_),
    .X(_2257_));
 sky130_fd_sc_hd__buf_1 _5028_ (.A(_2257_),
    .X(_0323_));
 sky130_fd_sc_hd__mux2_2 _5029_ (.A0(\tree_instances[14].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[14].u_tree.pipeline_frame_id[0][2] ),
    .S(_0735_),
    .X(_2258_));
 sky130_fd_sc_hd__buf_1 _5030_ (.A(_2258_),
    .X(_0324_));
 sky130_fd_sc_hd__mux2_2 _5031_ (.A0(\tree_instances[14].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[14].u_tree.pipeline_frame_id[0][3] ),
    .S(_0735_),
    .X(_2259_));
 sky130_fd_sc_hd__buf_1 _5032_ (.A(_2259_),
    .X(_0325_));
 sky130_fd_sc_hd__mux2_2 _5033_ (.A0(\tree_instances[14].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[14].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[14].u_tree.tree_state[3] ),
    .X(_2260_));
 sky130_fd_sc_hd__buf_1 _5034_ (.A(_2260_),
    .X(_0326_));
 sky130_fd_sc_hd__and2_2 _5035_ (.A(_1666_),
    .B(_2222_),
    .X(_2261_));
 sky130_fd_sc_hd__buf_1 _5036_ (.A(_2261_),
    .X(_0327_));
 sky130_fd_sc_hd__and2_2 _5037_ (.A(_1679_),
    .B(_2222_),
    .X(_2262_));
 sky130_fd_sc_hd__buf_1 _5038_ (.A(_2262_),
    .X(_0328_));
 sky130_fd_sc_hd__and2_2 _5039_ (.A(_1686_),
    .B(_2222_),
    .X(_2263_));
 sky130_fd_sc_hd__buf_1 _5040_ (.A(_2263_),
    .X(_0329_));
 sky130_fd_sc_hd__and2_2 _5041_ (.A(_1684_),
    .B(_2222_),
    .X(_2264_));
 sky130_fd_sc_hd__buf_1 _5042_ (.A(_2264_),
    .X(_0330_));
 sky130_fd_sc_hd__and2_2 _5043_ (.A(_1647_),
    .B(_2222_),
    .X(_2265_));
 sky130_fd_sc_hd__buf_1 _5044_ (.A(_2265_),
    .X(_0331_));
 sky130_fd_sc_hd__and2_2 _5045_ (.A(_1676_),
    .B(_2222_),
    .X(_2266_));
 sky130_fd_sc_hd__buf_1 _5046_ (.A(_2266_),
    .X(_0332_));
 sky130_fd_sc_hd__and2_2 _5047_ (.A(_1669_),
    .B(_2222_),
    .X(_2267_));
 sky130_fd_sc_hd__buf_1 _5048_ (.A(_2267_),
    .X(_0333_));
 sky130_fd_sc_hd__and2_2 _5049_ (.A(_1673_),
    .B(_2221_),
    .X(_2268_));
 sky130_fd_sc_hd__buf_1 _5050_ (.A(_2268_),
    .X(_0334_));
 sky130_fd_sc_hd__nand2_2 _5051_ (.A(\tree_instances[14].u_tree.tree_state[0] ),
    .B(_0734_),
    .Y(_2269_));
 sky130_fd_sc_hd__a22o_2 _5052_ (.A1(_0735_),
    .A2(_2269_),
    .B1(_1817_),
    .B2(\tree_instances[14].u_tree.ready_for_next ),
    .X(_0335_));
 sky130_fd_sc_hd__mux2_2 _5053_ (.A0(\tree_instances[15].u_tree.pipeline_frame_id[0][0] ),
    .A1(_2122_),
    .S(_0016_),
    .X(_2270_));
 sky130_fd_sc_hd__buf_1 _5054_ (.A(_2270_),
    .X(_0336_));
 sky130_fd_sc_hd__mux2_2 _5055_ (.A0(\tree_instances[15].u_tree.pipeline_frame_id[0][1] ),
    .A1(_2246_),
    .S(_0016_),
    .X(_2271_));
 sky130_fd_sc_hd__buf_1 _5056_ (.A(_2271_),
    .X(_0337_));
 sky130_fd_sc_hd__mux2_2 _5057_ (.A0(\tree_instances[15].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2125_),
    .S(_0016_),
    .X(_2272_));
 sky130_fd_sc_hd__buf_1 _5058_ (.A(_2272_),
    .X(_0338_));
 sky130_fd_sc_hd__mux2_2 _5059_ (.A0(\tree_instances[15].u_tree.pipeline_frame_id[0][3] ),
    .A1(_2249_),
    .S(_0016_),
    .X(_2273_));
 sky130_fd_sc_hd__buf_1 _5060_ (.A(_2273_),
    .X(_0339_));
 sky130_fd_sc_hd__mux2_2 _5061_ (.A0(\tree_instances[15].u_tree.pipeline_frame_id[0][4] ),
    .A1(_2251_),
    .S(_0016_),
    .X(_2274_));
 sky130_fd_sc_hd__buf_1 _5062_ (.A(_2274_),
    .X(_0340_));
 sky130_fd_sc_hd__inv_2 _5063_ (.A(_0016_),
    .Y(_2275_));
 sky130_fd_sc_hd__mux2_2 _5064_ (.A0(\tree_instances[15].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[15].u_tree.pipeline_frame_id[0][0] ),
    .S(_1137_),
    .X(_2276_));
 sky130_fd_sc_hd__buf_1 _5065_ (.A(_2276_),
    .X(_0341_));
 sky130_fd_sc_hd__mux2_2 _5066_ (.A0(\tree_instances[15].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[15].u_tree.pipeline_frame_id[0][1] ),
    .S(_1137_),
    .X(_2277_));
 sky130_fd_sc_hd__buf_1 _5067_ (.A(_2277_),
    .X(_0342_));
 sky130_fd_sc_hd__mux2_2 _5068_ (.A0(\tree_instances[15].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[15].u_tree.pipeline_frame_id[0][2] ),
    .S(_1137_),
    .X(_2278_));
 sky130_fd_sc_hd__buf_1 _5069_ (.A(_2278_),
    .X(_0343_));
 sky130_fd_sc_hd__mux2_2 _5070_ (.A0(\tree_instances[15].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[15].u_tree.pipeline_frame_id[0][3] ),
    .S(_1137_),
    .X(_2279_));
 sky130_fd_sc_hd__buf_1 _5071_ (.A(_2279_),
    .X(_0344_));
 sky130_fd_sc_hd__mux2_2 _5072_ (.A0(\tree_instances[15].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[15].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[15].u_tree.tree_state[3] ),
    .X(_2280_));
 sky130_fd_sc_hd__buf_1 _5073_ (.A(_2280_),
    .X(_0345_));
 sky130_fd_sc_hd__and2_2 _5074_ (.A(_1534_),
    .B(_2255_),
    .X(_2281_));
 sky130_fd_sc_hd__buf_1 _5075_ (.A(_2281_),
    .X(_0346_));
 sky130_fd_sc_hd__and2_2 _5076_ (.A(_1546_),
    .B(_2255_),
    .X(_2282_));
 sky130_fd_sc_hd__buf_1 _5077_ (.A(_2282_),
    .X(_0347_));
 sky130_fd_sc_hd__and2_2 _5078_ (.A(_1542_),
    .B(_2255_),
    .X(_2283_));
 sky130_fd_sc_hd__buf_1 _5079_ (.A(_2283_),
    .X(_0348_));
 sky130_fd_sc_hd__and2_2 _5080_ (.A(_1544_),
    .B(_2255_),
    .X(_2284_));
 sky130_fd_sc_hd__buf_1 _5081_ (.A(_2284_),
    .X(_0349_));
 sky130_fd_sc_hd__and2_2 _5082_ (.A(_1547_),
    .B(_2255_),
    .X(_2285_));
 sky130_fd_sc_hd__buf_1 _5083_ (.A(_2285_),
    .X(_0350_));
 sky130_fd_sc_hd__and2_2 _5084_ (.A(_1543_),
    .B(_2255_),
    .X(_2286_));
 sky130_fd_sc_hd__buf_1 _5085_ (.A(_2286_),
    .X(_0351_));
 sky130_fd_sc_hd__and2_2 _5086_ (.A(_1082_),
    .B(_2255_),
    .X(_2287_));
 sky130_fd_sc_hd__buf_1 _5087_ (.A(_2287_),
    .X(_0352_));
 sky130_fd_sc_hd__and2_2 _5088_ (.A(_1083_),
    .B(_2254_),
    .X(_2288_));
 sky130_fd_sc_hd__buf_1 _5089_ (.A(_2288_),
    .X(_0353_));
 sky130_fd_sc_hd__inv_2 _5090_ (.A(_1138_),
    .Y(_2289_));
 sky130_fd_sc_hd__a22o_2 _5091_ (.A1(_1137_),
    .A2(_2289_),
    .B1(_2275_),
    .B2(\tree_instances[15].u_tree.ready_for_next ),
    .X(_0354_));
 sky130_fd_sc_hd__buf_1 _5092_ (.A(\tree_instances[16].u_tree.tree_state[2] ),
    .X(_2290_));
 sky130_fd_sc_hd__a22o_2 _5093_ (.A1(\tree_instances[16].u_tree.tree_state[1] ),
    .A2(\tree_instances[16].u_tree.current_node_data[12] ),
    .B1(\tree_instances[16].u_tree.node_data[12] ),
    .B2(_2290_),
    .X(_2291_));
 sky130_fd_sc_hd__nor3_2 _5094_ (.A(\tree_instances[16].u_tree.tree_state[1] ),
    .B(\tree_instances[16].u_tree.tree_state[2] ),
    .C(\tree_instances[16].u_tree.tree_state[0] ),
    .Y(_2292_));
 sky130_fd_sc_hd__a211oi_2 _5095_ (.A1(\tree_instances[16].u_tree.tree_state[0] ),
    .A2(_1022_),
    .B1(_0017_),
    .C1(_2292_),
    .Y(_2293_));
 sky130_fd_sc_hd__mux2_2 _5096_ (.A0(\tree_instances[16].u_tree.pipeline_prediction[0][0] ),
    .A1(_2291_),
    .S(_2293_),
    .X(_2294_));
 sky130_fd_sc_hd__buf_1 _5097_ (.A(_2294_),
    .X(_0355_));
 sky130_fd_sc_hd__or2_2 _5098_ (.A(\tree_instances[16].u_tree.u_tree_weight_rom.cache_valid ),
    .B(\tree_instances[16].u_tree.read_enable ),
    .X(_2295_));
 sky130_fd_sc_hd__buf_1 _5099_ (.A(_2295_),
    .X(_0356_));
 sky130_fd_sc_hd__or3_2 _5100_ (.A(\tree_instances[15].u_tree.tree_state[2] ),
    .B(\tree_instances[15].u_tree.tree_state[1] ),
    .C(_2275_),
    .X(_2296_));
 sky130_fd_sc_hd__and2_2 _5101_ (.A(_1442_),
    .B(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__buf_1 _5102_ (.A(_2297_),
    .X(_0357_));
 sky130_fd_sc_hd__and2_2 _5103_ (.A(_1455_),
    .B(_2296_),
    .X(_2298_));
 sky130_fd_sc_hd__buf_1 _5104_ (.A(_2298_),
    .X(_0358_));
 sky130_fd_sc_hd__and2_2 _5105_ (.A(_1454_),
    .B(_2296_),
    .X(_2299_));
 sky130_fd_sc_hd__buf_1 _5106_ (.A(_2299_),
    .X(_0359_));
 sky130_fd_sc_hd__and2_2 _5107_ (.A(_1457_),
    .B(_2296_),
    .X(_2300_));
 sky130_fd_sc_hd__buf_1 _5108_ (.A(_2300_),
    .X(_0360_));
 sky130_fd_sc_hd__and2_2 _5109_ (.A(_1456_),
    .B(_2296_),
    .X(_2301_));
 sky130_fd_sc_hd__buf_1 _5110_ (.A(_2301_),
    .X(_0361_));
 sky130_fd_sc_hd__and2_2 _5111_ (.A(_1453_),
    .B(_2296_),
    .X(_2302_));
 sky130_fd_sc_hd__buf_1 _5112_ (.A(_2302_),
    .X(_0362_));
 sky130_fd_sc_hd__and2_2 _5113_ (.A(_1451_),
    .B(_2296_),
    .X(_2303_));
 sky130_fd_sc_hd__buf_1 _5114_ (.A(_2303_),
    .X(_0363_));
 sky130_fd_sc_hd__and2_2 _5115_ (.A(_1444_),
    .B(_2296_),
    .X(_2304_));
 sky130_fd_sc_hd__buf_1 _5116_ (.A(_2304_),
    .X(_0364_));
 sky130_fd_sc_hd__mux2_2 _5117_ (.A0(\tree_instances[16].u_tree.pipeline_frame_id[0][0] ),
    .A1(_2122_),
    .S(_0018_),
    .X(_2305_));
 sky130_fd_sc_hd__buf_1 _5118_ (.A(_2305_),
    .X(_0365_));
 sky130_fd_sc_hd__mux2_2 _5119_ (.A0(\tree_instances[16].u_tree.pipeline_frame_id[0][1] ),
    .A1(_2246_),
    .S(_0018_),
    .X(_2306_));
 sky130_fd_sc_hd__buf_1 _5120_ (.A(_2306_),
    .X(_0366_));
 sky130_fd_sc_hd__mux2_2 _5121_ (.A0(\tree_instances[16].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2125_),
    .S(_0018_),
    .X(_2307_));
 sky130_fd_sc_hd__buf_1 _5122_ (.A(_2307_),
    .X(_0367_));
 sky130_fd_sc_hd__mux2_2 _5123_ (.A0(\tree_instances[16].u_tree.pipeline_frame_id[0][3] ),
    .A1(_2249_),
    .S(_0018_),
    .X(_2308_));
 sky130_fd_sc_hd__buf_1 _5124_ (.A(_2308_),
    .X(_0368_));
 sky130_fd_sc_hd__mux2_2 _5125_ (.A0(\tree_instances[16].u_tree.pipeline_frame_id[0][4] ),
    .A1(_2251_),
    .S(_0018_),
    .X(_2309_));
 sky130_fd_sc_hd__buf_1 _5126_ (.A(_2309_),
    .X(_0369_));
 sky130_fd_sc_hd__inv_2 _5127_ (.A(\tree_instances[16].u_tree.read_enable ),
    .Y(_2310_));
 sky130_fd_sc_hd__buf_1 _5128_ (.A(_2310_),
    .X(_2311_));
 sky130_fd_sc_hd__nor2_2 _5129_ (.A(\tree_instances[16].u_tree.tree_state[1] ),
    .B(_2292_),
    .Y(_2312_));
 sky130_fd_sc_hd__or3_2 _5130_ (.A(\tree_instances[16].u_tree.tree_state[1] ),
    .B(\tree_instances[16].u_tree.tree_state[2] ),
    .C(_1809_),
    .X(_2313_));
 sky130_fd_sc_hd__buf_1 _5131_ (.A(_2313_),
    .X(_2314_));
 sky130_fd_sc_hd__o21ai_2 _5132_ (.A1(_2311_),
    .A2(_2312_),
    .B1(_2314_),
    .Y(_0370_));
 sky130_fd_sc_hd__mux2_2 _5133_ (.A0(\tree_instances[16].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[16].u_tree.pipeline_frame_id[0][0] ),
    .S(_1023_),
    .X(_2315_));
 sky130_fd_sc_hd__buf_1 _5134_ (.A(_2315_),
    .X(_0371_));
 sky130_fd_sc_hd__mux2_2 _5135_ (.A0(\tree_instances[16].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[16].u_tree.pipeline_frame_id[0][1] ),
    .S(_1023_),
    .X(_2316_));
 sky130_fd_sc_hd__buf_1 _5136_ (.A(_2316_),
    .X(_0372_));
 sky130_fd_sc_hd__mux2_2 _5137_ (.A0(\tree_instances[16].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[16].u_tree.pipeline_frame_id[0][2] ),
    .S(_1023_),
    .X(_2317_));
 sky130_fd_sc_hd__buf_1 _5138_ (.A(_2317_),
    .X(_0373_));
 sky130_fd_sc_hd__mux2_2 _5139_ (.A0(\tree_instances[16].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[16].u_tree.pipeline_frame_id[0][3] ),
    .S(_1023_),
    .X(_2318_));
 sky130_fd_sc_hd__buf_1 _5140_ (.A(_2318_),
    .X(_0374_));
 sky130_fd_sc_hd__mux2_2 _5141_ (.A0(\tree_instances[16].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[16].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[16].u_tree.tree_state[3] ),
    .X(_2319_));
 sky130_fd_sc_hd__buf_1 _5142_ (.A(_2319_),
    .X(_0375_));
 sky130_fd_sc_hd__mux2_2 _5143_ (.A0(\tree_instances[16].u_tree.prediction_out ),
    .A1(\tree_instances[16].u_tree.pipeline_prediction[0][0] ),
    .S(\tree_instances[16].u_tree.tree_state[3] ),
    .X(_2320_));
 sky130_fd_sc_hd__buf_1 _5144_ (.A(_2320_),
    .X(_0376_));
 sky130_fd_sc_hd__nand2_2 _5145_ (.A(\tree_instances[16].u_tree.tree_state[0] ),
    .B(_1022_),
    .Y(_2321_));
 sky130_fd_sc_hd__a22o_2 _5146_ (.A1(_1023_),
    .A2(_2321_),
    .B1(_1809_),
    .B2(\tree_instances[16].u_tree.ready_for_next ),
    .X(_0377_));
 sky130_fd_sc_hd__nand2_2 _5147_ (.A(\tree_instances[14].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[14].u_tree.tree_state[0] ),
    .Y(_2322_));
 sky130_fd_sc_hd__o2bb2a_2 _5148_ (.A1_N(_0735_),
    .A2_N(_2322_),
    .B1(_0014_),
    .B2(\tree_instances[14].u_tree.pipeline_valid[0] ),
    .X(_0378_));
 sky130_fd_sc_hd__buf_1 _5149_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][3] ),
    .X(_2323_));
 sky130_fd_sc_hd__buf_1 _5150_ (.A(_0786_),
    .X(_2324_));
 sky130_fd_sc_hd__buf_1 _5151_ (.A(_2324_),
    .X(_2325_));
 sky130_fd_sc_hd__buf_1 _5152_ (.A(_0785_),
    .X(_2326_));
 sky130_fd_sc_hd__buf_1 _5153_ (.A(_0781_),
    .X(_2327_));
 sky130_fd_sc_hd__buf_1 _5154_ (.A(_2327_),
    .X(_2328_));
 sky130_fd_sc_hd__buf_1 _5155_ (.A(_2323_),
    .X(_2329_));
 sky130_fd_sc_hd__buf_1 _5156_ (.A(_2329_),
    .X(_2330_));
 sky130_fd_sc_hd__buf_1 _5157_ (.A(_2330_),
    .X(_2331_));
 sky130_fd_sc_hd__buf_1 _5158_ (.A(_2331_),
    .X(_2332_));
 sky130_fd_sc_hd__buf_1 _5159_ (.A(_0793_),
    .X(_2333_));
 sky130_fd_sc_hd__buf_1 _5160_ (.A(_2333_),
    .X(_2334_));
 sky130_fd_sc_hd__buf_1 _5161_ (.A(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__buf_1 _5162_ (.A(_2335_),
    .X(_2336_));
 sky130_fd_sc_hd__buf_1 _5163_ (.A(_0792_),
    .X(_2337_));
 sky130_fd_sc_hd__buf_1 _5164_ (.A(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__buf_1 _5165_ (.A(_2338_),
    .X(_2339_));
 sky130_fd_sc_hd__buf_1 _5166_ (.A(_2339_),
    .X(_2340_));
 sky130_fd_sc_hd__buf_1 _5167_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][6] ),
    .X(_2341_));
 sky130_fd_sc_hd__buf_1 _5168_ (.A(_2341_),
    .X(_2342_));
 sky130_fd_sc_hd__buf_1 _5169_ (.A(_2342_),
    .X(_2343_));
 sky130_fd_sc_hd__buf_1 _5170_ (.A(_2343_),
    .X(_2344_));
 sky130_fd_sc_hd__buf_1 _5171_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][7] ),
    .X(_2345_));
 sky130_fd_sc_hd__buf_1 _5172_ (.A(_2345_),
    .X(_2346_));
 sky130_fd_sc_hd__inv_2 _5173_ (.A(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .Y(_2347_));
 sky130_fd_sc_hd__inv_2 _5174_ (.A(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .Y(_2348_));
 sky130_fd_sc_hd__nor2_2 _5175_ (.A(_1371_),
    .B(_2348_),
    .Y(_2349_));
 sky130_fd_sc_hd__a221o_2 _5176_ (.A1(\tree_instances[16].u_tree.pipeline_current_node[0][6] ),
    .A2(_2347_),
    .B1(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .B2(_1368_),
    .C1(_2349_),
    .X(_2350_));
 sky130_fd_sc_hd__xor2_2 _5177_ (.A(_1367_),
    .B(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .X(_2351_));
 sky130_fd_sc_hd__a221o_2 _5178_ (.A1(_1375_),
    .A2(_2348_),
    .B1(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .B2(_1355_),
    .C1(_2351_),
    .X(_2352_));
 sky130_fd_sc_hd__nor2_2 _5179_ (.A(_1217_),
    .B(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .Y(_2353_));
 sky130_fd_sc_hd__and2_2 _5180_ (.A(_1217_),
    .B(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .X(_2354_));
 sky130_fd_sc_hd__xnor2_2 _5181_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][5] ),
    .B(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .Y(_2355_));
 sky130_fd_sc_hd__o221a_2 _5182_ (.A1(_1355_),
    .A2(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .B1(_2353_),
    .B2(_2354_),
    .C1(_2355_),
    .X(_2356_));
 sky130_fd_sc_hd__xnor2_2 _5183_ (.A(\tree_instances[16].u_tree.pipeline_current_node[0][4] ),
    .B(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .Y(_2357_));
 sky130_fd_sc_hd__o221a_2 _5184_ (.A1(\tree_instances[16].u_tree.pipeline_current_node[0][6] ),
    .A2(_2347_),
    .B1(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .B2(_1368_),
    .C1(_2357_),
    .X(_2358_));
 sky130_fd_sc_hd__and3_2 _5185_ (.A(\tree_instances[16].u_tree.u_tree_weight_rom.cache_valid ),
    .B(_2356_),
    .C(_2358_),
    .X(_2359_));
 sky130_fd_sc_hd__or3b_2 _5186_ (.A(_2350_),
    .B(_2352_),
    .C_N(_2359_),
    .X(_2360_));
 sky130_fd_sc_hd__and2_2 _5187_ (.A(\tree_instances[16].u_tree.read_enable ),
    .B(_2360_),
    .X(_2361_));
 sky130_fd_sc_hd__buf_1 _5188_ (.A(_2361_),
    .X(_2362_));
 sky130_fd_sc_hd__buf_1 _5189_ (.A(_2362_),
    .X(_2363_));
 sky130_fd_sc_hd__mux2_2 _5190_ (.A0(\tree_instances[16].u_tree.u_tree_weight_rom.cached_data[12] ),
    .A1(\tree_instances[16].u_tree.u_tree_weight_rom.gen_tree_16.u_tree_rom.node_data[12] ),
    .S(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__buf_1 _5191_ (.A(_2364_),
    .X(_0380_));
 sky130_fd_sc_hd__inv_2 _5192_ (.A(_0020_),
    .Y(_2365_));
 sky130_fd_sc_hd__or3_2 _5193_ (.A(\tree_instances[17].u_tree.tree_state[2] ),
    .B(\tree_instances[17].u_tree.tree_state[1] ),
    .C(_2365_),
    .X(_2366_));
 sky130_fd_sc_hd__buf_1 _5194_ (.A(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__and2_2 _5195_ (.A(_2325_),
    .B(_2367_),
    .X(_2368_));
 sky130_fd_sc_hd__buf_1 _5196_ (.A(_2368_),
    .X(_0381_));
 sky130_fd_sc_hd__and2_2 _5197_ (.A(_2326_),
    .B(_2367_),
    .X(_2369_));
 sky130_fd_sc_hd__buf_1 _5198_ (.A(_2369_),
    .X(_0382_));
 sky130_fd_sc_hd__and2_2 _5199_ (.A(_2328_),
    .B(_2367_),
    .X(_2370_));
 sky130_fd_sc_hd__buf_1 _5200_ (.A(_2370_),
    .X(_0383_));
 sky130_fd_sc_hd__and2_2 _5201_ (.A(_2332_),
    .B(_2367_),
    .X(_2371_));
 sky130_fd_sc_hd__buf_1 _5202_ (.A(_2371_),
    .X(_0384_));
 sky130_fd_sc_hd__and2_2 _5203_ (.A(_2336_),
    .B(_2367_),
    .X(_2372_));
 sky130_fd_sc_hd__buf_1 _5204_ (.A(_2372_),
    .X(_0385_));
 sky130_fd_sc_hd__and2_2 _5205_ (.A(_2340_),
    .B(_2367_),
    .X(_2373_));
 sky130_fd_sc_hd__buf_1 _5206_ (.A(_2373_),
    .X(_0386_));
 sky130_fd_sc_hd__and2_2 _5207_ (.A(_2344_),
    .B(_2367_),
    .X(_2374_));
 sky130_fd_sc_hd__buf_1 _5208_ (.A(_2374_),
    .X(_0387_));
 sky130_fd_sc_hd__and2_2 _5209_ (.A(_2346_),
    .B(_2367_),
    .X(_2375_));
 sky130_fd_sc_hd__buf_1 _5210_ (.A(_2375_),
    .X(_0388_));
 sky130_fd_sc_hd__buf_1 _5211_ (.A(\tree_instances[17].u_tree.pipeline_current_node[0][8] ),
    .X(_2376_));
 sky130_fd_sc_hd__and2_2 _5212_ (.A(_2376_),
    .B(_2366_),
    .X(_2377_));
 sky130_fd_sc_hd__buf_1 _5213_ (.A(_2377_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_2 _5214_ (.A0(\tree_instances[17].u_tree.pipeline_frame_id[0][0] ),
    .A1(_2122_),
    .S(_0020_),
    .X(_2378_));
 sky130_fd_sc_hd__buf_1 _5215_ (.A(_2378_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_2 _5216_ (.A0(\tree_instances[17].u_tree.pipeline_frame_id[0][1] ),
    .A1(_2246_),
    .S(_0020_),
    .X(_2379_));
 sky130_fd_sc_hd__buf_1 _5217_ (.A(_2379_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_2 _5218_ (.A0(\tree_instances[17].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2125_),
    .S(_0020_),
    .X(_2380_));
 sky130_fd_sc_hd__buf_1 _5219_ (.A(_2380_),
    .X(_0392_));
 sky130_fd_sc_hd__mux2_2 _5220_ (.A0(\tree_instances[17].u_tree.pipeline_frame_id[0][3] ),
    .A1(_2249_),
    .S(_0020_),
    .X(_2381_));
 sky130_fd_sc_hd__buf_1 _5221_ (.A(_2381_),
    .X(_0393_));
 sky130_fd_sc_hd__mux2_2 _5222_ (.A0(\tree_instances[17].u_tree.pipeline_frame_id[0][4] ),
    .A1(_2251_),
    .S(_0020_),
    .X(_2382_));
 sky130_fd_sc_hd__buf_1 _5223_ (.A(_2382_),
    .X(_0394_));
 sky130_fd_sc_hd__mux2_2 _5224_ (.A0(\tree_instances[16].u_tree.current_node_data[12] ),
    .A1(\tree_instances[16].u_tree.node_data[12] ),
    .S(_0912_),
    .X(_2383_));
 sky130_fd_sc_hd__buf_1 _5225_ (.A(_2383_),
    .X(_0395_));
 sky130_fd_sc_hd__mux2_2 _5226_ (.A0(\tree_instances[17].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[17].u_tree.pipeline_frame_id[0][0] ),
    .S(_0909_),
    .X(_2384_));
 sky130_fd_sc_hd__buf_1 _5227_ (.A(_2384_),
    .X(_0396_));
 sky130_fd_sc_hd__mux2_2 _5228_ (.A0(\tree_instances[17].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[17].u_tree.pipeline_frame_id[0][1] ),
    .S(_0909_),
    .X(_2385_));
 sky130_fd_sc_hd__buf_1 _5229_ (.A(_2385_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_2 _5230_ (.A0(\tree_instances[17].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[17].u_tree.pipeline_frame_id[0][2] ),
    .S(_0909_),
    .X(_2386_));
 sky130_fd_sc_hd__buf_1 _5231_ (.A(_2386_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_2 _5232_ (.A0(\tree_instances[17].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[17].u_tree.pipeline_frame_id[0][3] ),
    .S(_0909_),
    .X(_2387_));
 sky130_fd_sc_hd__buf_1 _5233_ (.A(_2387_),
    .X(_0399_));
 sky130_fd_sc_hd__mux2_2 _5234_ (.A0(\tree_instances[17].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[17].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[17].u_tree.tree_state[3] ),
    .X(_2388_));
 sky130_fd_sc_hd__buf_1 _5235_ (.A(_2388_),
    .X(_0400_));
 sky130_fd_sc_hd__and2_2 _5236_ (.A(_1386_),
    .B(_2314_),
    .X(_2389_));
 sky130_fd_sc_hd__buf_1 _5237_ (.A(_2389_),
    .X(_0401_));
 sky130_fd_sc_hd__and2_2 _5238_ (.A(_1379_),
    .B(_2314_),
    .X(_2390_));
 sky130_fd_sc_hd__buf_1 _5239_ (.A(_2390_),
    .X(_0402_));
 sky130_fd_sc_hd__and2_2 _5240_ (.A(_1382_),
    .B(_2314_),
    .X(_2391_));
 sky130_fd_sc_hd__buf_1 _5241_ (.A(_2391_),
    .X(_0403_));
 sky130_fd_sc_hd__and2_2 _5242_ (.A(_1384_),
    .B(_2314_),
    .X(_2392_));
 sky130_fd_sc_hd__buf_1 _5243_ (.A(_2392_),
    .X(_0404_));
 sky130_fd_sc_hd__and2_2 _5244_ (.A(_1380_),
    .B(_2314_),
    .X(_2393_));
 sky130_fd_sc_hd__buf_1 _5245_ (.A(_2393_),
    .X(_0405_));
 sky130_fd_sc_hd__and2_2 _5246_ (.A(_1383_),
    .B(_2314_),
    .X(_2394_));
 sky130_fd_sc_hd__buf_1 _5247_ (.A(_2394_),
    .X(_0406_));
 sky130_fd_sc_hd__and2_2 _5248_ (.A(_1388_),
    .B(_2314_),
    .X(_2395_));
 sky130_fd_sc_hd__buf_1 _5249_ (.A(_2395_),
    .X(_0407_));
 sky130_fd_sc_hd__and2_2 _5250_ (.A(_1385_),
    .B(_2313_),
    .X(_2396_));
 sky130_fd_sc_hd__buf_1 _5251_ (.A(_2396_),
    .X(_0408_));
 sky130_fd_sc_hd__inv_2 _5252_ (.A(_0910_),
    .Y(_2397_));
 sky130_fd_sc_hd__a22o_2 _5253_ (.A1(_0909_),
    .A2(_2397_),
    .B1(_2365_),
    .B2(\tree_instances[17].u_tree.ready_for_next ),
    .X(_0409_));
 sky130_fd_sc_hd__nand2_2 _5254_ (.A(\tree_instances[9].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[9].u_tree.tree_state[0] ),
    .Y(_2398_));
 sky130_fd_sc_hd__o2bb2a_2 _5255_ (.A1_N(_1025_),
    .A2_N(_2398_),
    .B1(_0044_),
    .B2(\tree_instances[9].u_tree.pipeline_valid[0] ),
    .X(_0410_));
 sky130_fd_sc_hd__buf_1 _5256_ (.A(_2362_),
    .X(_2399_));
 sky130_fd_sc_hd__mux2_2 _5257_ (.A0(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .A1(_1386_),
    .S(_2399_),
    .X(_2400_));
 sky130_fd_sc_hd__buf_1 _5258_ (.A(_2400_),
    .X(_0411_));
 sky130_fd_sc_hd__mux2_2 _5259_ (.A0(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .A1(_1379_),
    .S(_2399_),
    .X(_2401_));
 sky130_fd_sc_hd__buf_1 _5260_ (.A(_2401_),
    .X(_0412_));
 sky130_fd_sc_hd__mux2_2 _5261_ (.A0(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .A1(_1382_),
    .S(_2399_),
    .X(_2402_));
 sky130_fd_sc_hd__buf_1 _5262_ (.A(_2402_),
    .X(_0413_));
 sky130_fd_sc_hd__mux2_2 _5263_ (.A0(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .A1(_1384_),
    .S(_2399_),
    .X(_2403_));
 sky130_fd_sc_hd__buf_1 _5264_ (.A(_2403_),
    .X(_0414_));
 sky130_fd_sc_hd__mux2_2 _5265_ (.A0(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .A1(_1380_),
    .S(_2399_),
    .X(_2404_));
 sky130_fd_sc_hd__buf_1 _5266_ (.A(_2404_),
    .X(_0415_));
 sky130_fd_sc_hd__mux2_2 _5267_ (.A0(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .A1(_1383_),
    .S(_2399_),
    .X(_2405_));
 sky130_fd_sc_hd__buf_1 _5268_ (.A(_2405_),
    .X(_0416_));
 sky130_fd_sc_hd__mux2_2 _5269_ (.A0(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .A1(_1388_),
    .S(_2399_),
    .X(_2406_));
 sky130_fd_sc_hd__buf_1 _5270_ (.A(_2406_),
    .X(_0417_));
 sky130_fd_sc_hd__mux2_2 _5271_ (.A0(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .A1(_1376_),
    .S(_2399_),
    .X(_2407_));
 sky130_fd_sc_hd__buf_1 _5272_ (.A(_2407_),
    .X(_0418_));
 sky130_fd_sc_hd__mux2_2 _5273_ (.A0(\tree_instances[18].u_tree.pipeline_frame_id[0][0] ),
    .A1(_2122_),
    .S(_0022_),
    .X(_2408_));
 sky130_fd_sc_hd__buf_1 _5274_ (.A(_2408_),
    .X(_0419_));
 sky130_fd_sc_hd__mux2_2 _5275_ (.A0(\tree_instances[18].u_tree.pipeline_frame_id[0][1] ),
    .A1(_2246_),
    .S(_0022_),
    .X(_2409_));
 sky130_fd_sc_hd__buf_1 _5276_ (.A(_2409_),
    .X(_0420_));
 sky130_fd_sc_hd__mux2_2 _5277_ (.A0(\tree_instances[18].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2125_),
    .S(_0022_),
    .X(_2410_));
 sky130_fd_sc_hd__buf_1 _5278_ (.A(_2410_),
    .X(_0421_));
 sky130_fd_sc_hd__mux2_2 _5279_ (.A0(\tree_instances[18].u_tree.pipeline_frame_id[0][3] ),
    .A1(_2249_),
    .S(_0022_),
    .X(_2411_));
 sky130_fd_sc_hd__buf_1 _5280_ (.A(_2411_),
    .X(_0422_));
 sky130_fd_sc_hd__mux2_2 _5281_ (.A0(\tree_instances[18].u_tree.pipeline_frame_id[0][4] ),
    .A1(_2251_),
    .S(_0022_),
    .X(_2412_));
 sky130_fd_sc_hd__buf_1 _5282_ (.A(_2412_),
    .X(_0423_));
 sky130_fd_sc_hd__or3_2 _5283_ (.A(\tree_instances[18].u_tree.tree_state[1] ),
    .B(\tree_instances[18].u_tree.tree_state[2] ),
    .C(_1801_),
    .X(_2413_));
 sky130_fd_sc_hd__buf_1 _5284_ (.A(_2413_),
    .X(_2414_));
 sky130_fd_sc_hd__mux2_2 _5285_ (.A0(\tree_instances[18].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[18].u_tree.pipeline_frame_id[0][0] ),
    .S(_0753_),
    .X(_2415_));
 sky130_fd_sc_hd__buf_1 _5286_ (.A(_2415_),
    .X(_0424_));
 sky130_fd_sc_hd__mux2_2 _5287_ (.A0(\tree_instances[18].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[18].u_tree.pipeline_frame_id[0][1] ),
    .S(_0753_),
    .X(_2416_));
 sky130_fd_sc_hd__buf_1 _5288_ (.A(_2416_),
    .X(_0425_));
 sky130_fd_sc_hd__mux2_2 _5289_ (.A0(\tree_instances[18].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[18].u_tree.pipeline_frame_id[0][2] ),
    .S(_0753_),
    .X(_2417_));
 sky130_fd_sc_hd__buf_1 _5290_ (.A(_2417_),
    .X(_0426_));
 sky130_fd_sc_hd__mux2_2 _5291_ (.A0(\tree_instances[18].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[18].u_tree.pipeline_frame_id[0][3] ),
    .S(_0753_),
    .X(_2418_));
 sky130_fd_sc_hd__buf_1 _5292_ (.A(_2418_),
    .X(_0427_));
 sky130_fd_sc_hd__mux2_2 _5293_ (.A0(\tree_instances[18].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[18].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[18].u_tree.tree_state[3] ),
    .X(_2419_));
 sky130_fd_sc_hd__buf_1 _5294_ (.A(_2419_),
    .X(_0428_));
 sky130_fd_sc_hd__a22o_2 _5295_ (.A1(_0753_),
    .A2(_1884_),
    .B1(_1801_),
    .B2(\tree_instances[18].u_tree.ready_for_next ),
    .X(_0429_));
 sky130_fd_sc_hd__nand2_2 _5296_ (.A(\tree_instances[15].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[15].u_tree.tree_state[0] ),
    .Y(_2420_));
 sky130_fd_sc_hd__o2bb2a_2 _5297_ (.A1_N(_1137_),
    .A2_N(_2420_),
    .B1(_0016_),
    .B2(\tree_instances[15].u_tree.pipeline_valid[0] ),
    .X(_0430_));
 sky130_fd_sc_hd__mux2_2 _5298_ (.A0(\tree_instances[19].u_tree.pipeline_frame_id[0][0] ),
    .A1(_2122_),
    .S(_0024_),
    .X(_2421_));
 sky130_fd_sc_hd__buf_1 _5299_ (.A(_2421_),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_2 _5300_ (.A0(\tree_instances[19].u_tree.pipeline_frame_id[0][1] ),
    .A1(_2246_),
    .S(_0024_),
    .X(_2422_));
 sky130_fd_sc_hd__buf_1 _5301_ (.A(_2422_),
    .X(_0432_));
 sky130_fd_sc_hd__mux2_2 _5302_ (.A0(\tree_instances[19].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2125_),
    .S(_0024_),
    .X(_2423_));
 sky130_fd_sc_hd__buf_1 _5303_ (.A(_2423_),
    .X(_0433_));
 sky130_fd_sc_hd__mux2_2 _5304_ (.A0(\tree_instances[19].u_tree.pipeline_frame_id[0][3] ),
    .A1(_2249_),
    .S(_0024_),
    .X(_2424_));
 sky130_fd_sc_hd__buf_1 _5305_ (.A(_2424_),
    .X(_0434_));
 sky130_fd_sc_hd__mux2_2 _5306_ (.A0(\tree_instances[19].u_tree.pipeline_frame_id[0][4] ),
    .A1(_2251_),
    .S(_0024_),
    .X(_2425_));
 sky130_fd_sc_hd__buf_1 _5307_ (.A(_2425_),
    .X(_0435_));
 sky130_fd_sc_hd__or3_2 _5308_ (.A(\tree_instances[19].u_tree.tree_state[1] ),
    .B(\tree_instances[19].u_tree.tree_state[2] ),
    .C(_1825_),
    .X(_2426_));
 sky130_fd_sc_hd__buf_1 _5309_ (.A(_2426_),
    .X(_2427_));
 sky130_fd_sc_hd__mux2_2 _5310_ (.A0(\tree_instances[19].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[19].u_tree.pipeline_frame_id[0][0] ),
    .S(_1252_),
    .X(_2428_));
 sky130_fd_sc_hd__buf_1 _5311_ (.A(_2428_),
    .X(_0436_));
 sky130_fd_sc_hd__mux2_2 _5312_ (.A0(\tree_instances[19].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[19].u_tree.pipeline_frame_id[0][1] ),
    .S(_1252_),
    .X(_2429_));
 sky130_fd_sc_hd__buf_1 _5313_ (.A(_2429_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_2 _5314_ (.A0(\tree_instances[19].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[19].u_tree.pipeline_frame_id[0][2] ),
    .S(_1252_),
    .X(_2430_));
 sky130_fd_sc_hd__buf_1 _5315_ (.A(_2430_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_2 _5316_ (.A0(\tree_instances[19].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[19].u_tree.pipeline_frame_id[0][3] ),
    .S(_1252_),
    .X(_2431_));
 sky130_fd_sc_hd__buf_1 _5317_ (.A(_2431_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_2 _5318_ (.A0(\tree_instances[19].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[19].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[19].u_tree.tree_state[3] ),
    .X(_2432_));
 sky130_fd_sc_hd__buf_1 _5319_ (.A(_2432_),
    .X(_0440_));
 sky130_fd_sc_hd__and2_2 _5320_ (.A(_1568_),
    .B(_2414_),
    .X(_2433_));
 sky130_fd_sc_hd__buf_1 _5321_ (.A(_2433_),
    .X(_0441_));
 sky130_fd_sc_hd__and2_2 _5322_ (.A(_1571_),
    .B(_2414_),
    .X(_2434_));
 sky130_fd_sc_hd__buf_1 _5323_ (.A(_2434_),
    .X(_0442_));
 sky130_fd_sc_hd__and2_2 _5324_ (.A(_1572_),
    .B(_2414_),
    .X(_2435_));
 sky130_fd_sc_hd__buf_1 _5325_ (.A(_2435_),
    .X(_0443_));
 sky130_fd_sc_hd__and2_2 _5326_ (.A(_1566_),
    .B(_2414_),
    .X(_2436_));
 sky130_fd_sc_hd__buf_1 _5327_ (.A(_2436_),
    .X(_0444_));
 sky130_fd_sc_hd__and2_2 _5328_ (.A(_1570_),
    .B(_2414_),
    .X(_2437_));
 sky130_fd_sc_hd__buf_1 _5329_ (.A(_2437_),
    .X(_0445_));
 sky130_fd_sc_hd__and2_2 _5330_ (.A(_1569_),
    .B(_2414_),
    .X(_2438_));
 sky130_fd_sc_hd__buf_1 _5331_ (.A(_2438_),
    .X(_0446_));
 sky130_fd_sc_hd__and2_2 _5332_ (.A(_1564_),
    .B(_2414_),
    .X(_2439_));
 sky130_fd_sc_hd__buf_1 _5333_ (.A(_2439_),
    .X(_0447_));
 sky130_fd_sc_hd__and2_2 _5334_ (.A(_1561_),
    .B(_2413_),
    .X(_2440_));
 sky130_fd_sc_hd__buf_1 _5335_ (.A(_2440_),
    .X(_0448_));
 sky130_fd_sc_hd__a22o_2 _5336_ (.A1(_1252_),
    .A2(_1989_),
    .B1(_1825_),
    .B2(\tree_instances[19].u_tree.ready_for_next ),
    .X(_0449_));
 sky130_fd_sc_hd__or4_2 _5337_ (.A(_0731_),
    .B(_0993_),
    .C(_0996_),
    .D(_0998_),
    .X(_2441_));
 sky130_fd_sc_hd__or2b_2 _5338_ (.A(\state[0] ),
    .B_N(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__inv_2 _5339_ (.A(\complete_votes[4] ),
    .Y(_2443_));
 sky130_fd_sc_hd__nand2_2 _5340_ (.A(\complete_votes[0] ),
    .B(\complete_votes[2] ),
    .Y(_2444_));
 sky130_fd_sc_hd__or4_2 _5341_ (.A(\complete_votes[1] ),
    .B(\complete_votes[3] ),
    .C(_2443_),
    .D(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__and3_2 _5342_ (.A(_1018_),
    .B(_2442_),
    .C(_2445_),
    .X(_2446_));
 sky130_fd_sc_hd__buf_1 _5343_ (.A(_2446_),
    .X(_0450_));
 sky130_fd_sc_hd__buf_1 _5344_ (.A(\state[1] ),
    .X(_2447_));
 sky130_fd_sc_hd__nor2_2 _5345_ (.A(_2447_),
    .B(_2445_),
    .Y(_0451_));
 sky130_fd_sc_hd__buf_1 _5346_ (.A(_0938_),
    .X(_2448_));
 sky130_fd_sc_hd__buf_1 _5347_ (.A(_1240_),
    .X(_2449_));
 sky130_fd_sc_hd__inv_2 _5348_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][1] ),
    .Y(_2450_));
 sky130_fd_sc_hd__nor2_2 _5349_ (.A(_2449_),
    .B(_2450_),
    .Y(_2451_));
 sky130_fd_sc_hd__buf_1 _5350_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][3] ),
    .X(_2452_));
 sky130_fd_sc_hd__inv_2 _5351_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][4] ),
    .Y(_2453_));
 sky130_fd_sc_hd__buf_1 _5352_ (.A(_2453_),
    .X(_2454_));
 sky130_fd_sc_hd__buf_1 _5353_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][5] ),
    .X(_2455_));
 sky130_fd_sc_hd__buf_1 _5354_ (.A(_2449_),
    .X(_2456_));
 sky130_fd_sc_hd__nand2_2 _5355_ (.A(_2452_),
    .B(_0939_),
    .Y(_2457_));
 sky130_fd_sc_hd__buf_1 _5356_ (.A(_1248_),
    .X(_2458_));
 sky130_fd_sc_hd__inv_2 _5357_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][2] ),
    .Y(_2459_));
 sky130_fd_sc_hd__inv_2 _5358_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][0] ),
    .Y(_2460_));
 sky130_fd_sc_hd__buf_1 _5359_ (.A(_2455_),
    .X(_2461_));
 sky130_fd_sc_hd__buf_1 _5360_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][6] ),
    .X(_2462_));
 sky130_fd_sc_hd__buf_1 _5361_ (.A(_2462_),
    .X(_2463_));
 sky130_fd_sc_hd__inv_2 _5362_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][5] ),
    .Y(_2464_));
 sky130_fd_sc_hd__buf_1 _5363_ (.A(_2459_),
    .X(_2465_));
 sky130_fd_sc_hd__buf_1 _5364_ (.A(_2458_),
    .X(_2466_));
 sky130_fd_sc_hd__buf_1 _5365_ (.A(_2448_),
    .X(_2467_));
 sky130_fd_sc_hd__buf_1 _5366_ (.A(_2467_),
    .X(_2468_));
 sky130_fd_sc_hd__buf_1 _5367_ (.A(_2466_),
    .X(_2469_));
 sky130_fd_sc_hd__buf_1 _5368_ (.A(_0937_),
    .X(_2470_));
 sky130_fd_sc_hd__buf_1 _5369_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][1] ),
    .X(_2471_));
 sky130_fd_sc_hd__inv_2 _5370_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][8] ),
    .Y(_2472_));
 sky130_fd_sc_hd__buf_1 _5371_ (.A(_2472_),
    .X(_2473_));
 sky130_fd_sc_hd__buf_1 _5372_ (.A(_2463_),
    .X(_2474_));
 sky130_fd_sc_hd__buf_1 _5373_ (.A(_0944_),
    .X(_2475_));
 sky130_fd_sc_hd__buf_1 _5374_ (.A(_2461_),
    .X(_2476_));
 sky130_fd_sc_hd__buf_1 _5375_ (.A(_2476_),
    .X(_2477_));
 sky130_fd_sc_hd__buf_1 _5376_ (.A(_2465_),
    .X(_2478_));
 sky130_fd_sc_hd__nand2_2 _5377_ (.A(_1240_),
    .B(_2471_),
    .Y(_2479_));
 sky130_fd_sc_hd__buf_1 _5378_ (.A(_0940_),
    .X(_2480_));
 sky130_fd_sc_hd__buf_1 _5379_ (.A(_2480_),
    .X(_2481_));
 sky130_fd_sc_hd__buf_1 _5380_ (.A(_2479_),
    .X(_2482_));
 sky130_fd_sc_hd__and2_2 _5381_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][7] ),
    .B(_2473_),
    .X(_2483_));
 sky130_fd_sc_hd__buf_1 _5382_ (.A(_2483_),
    .X(_2484_));
 sky130_fd_sc_hd__nor2_2 _5383_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][5] ),
    .B(_1247_),
    .Y(_2485_));
 sky130_fd_sc_hd__buf_1 _5384_ (.A(_2471_),
    .X(_2486_));
 sky130_fd_sc_hd__nor2_2 _5385_ (.A(_2455_),
    .B(_2462_),
    .Y(_2487_));
 sky130_fd_sc_hd__nor2_2 _5386_ (.A(_2470_),
    .B(_2454_),
    .Y(_2488_));
 sky130_fd_sc_hd__nor2_2 _5387_ (.A(_2464_),
    .B(_1247_),
    .Y(_2489_));
 sky130_fd_sc_hd__buf_1 _5388_ (.A(_2469_),
    .X(_2490_));
 sky130_fd_sc_hd__buf_1 _5389_ (.A(_2487_),
    .X(_2491_));
 sky130_fd_sc_hd__nor2_2 _5390_ (.A(_2457_),
    .B(_2482_),
    .Y(_2492_));
 sky130_fd_sc_hd__and3_2 _5391_ (.A(_2491_),
    .B(_2451_),
    .C(_2488_),
    .X(_2493_));
 sky130_fd_sc_hd__nand2_2 _5392_ (.A(\tree_instances[8].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[8].u_tree.tree_state[0] ),
    .Y(_2494_));
 sky130_fd_sc_hd__o2bb2a_2 _5393_ (.A1_N(_1000_),
    .A2_N(_2494_),
    .B1(_0042_),
    .B2(\tree_instances[8].u_tree.pipeline_valid[0] ),
    .X(_0452_));
 sky130_fd_sc_hd__nand2_2 _5394_ (.A(\tree_instances[0].u_tree.tree_state[0] ),
    .B(_0736_),
    .Y(_2495_));
 sky130_fd_sc_hd__o2bb2a_2 _5395_ (.A1_N(_0737_),
    .A2_N(_2495_),
    .B1(_0004_),
    .B2(\tree_instances[0].u_tree.pipeline_valid[0] ),
    .X(_0453_));
 sky130_fd_sc_hd__nand2_2 _5396_ (.A(\tree_instances[10].u_tree.tree_state[0] ),
    .B(\tree_instances[10].u_tree.pipeline_valid[0] ),
    .Y(_2496_));
 sky130_fd_sc_hd__o2bb2a_2 _5397_ (.A1_N(_1136_),
    .A2_N(_2496_),
    .B1(_0006_),
    .B2(\tree_instances[10].u_tree.pipeline_valid[0] ),
    .X(_0454_));
 sky130_fd_sc_hd__buf_1 _5398_ (.A(_0756_),
    .X(_2497_));
 sky130_fd_sc_hd__a22o_2 _5399_ (.A1(\tree_instances[20].u_tree.tree_state[1] ),
    .A2(\tree_instances[20].u_tree.current_node_data[12] ),
    .B1(\tree_instances[20].u_tree.node_data[12] ),
    .B2(_2497_),
    .X(_2498_));
 sky130_fd_sc_hd__or3_2 _5400_ (.A(\tree_instances[20].u_tree.tree_state[2] ),
    .B(\tree_instances[20].u_tree.tree_state[1] ),
    .C(\tree_instances[20].u_tree.tree_state[0] ),
    .X(_2499_));
 sky130_fd_sc_hd__and3b_2 _5401_ (.A_N(_0027_),
    .B(_1198_),
    .C(_2499_),
    .X(_2500_));
 sky130_fd_sc_hd__mux2_2 _5402_ (.A0(\tree_instances[20].u_tree.pipeline_prediction[0][0] ),
    .A1(_2498_),
    .S(_2500_),
    .X(_2501_));
 sky130_fd_sc_hd__buf_1 _5403_ (.A(_2501_),
    .X(_0455_));
 sky130_fd_sc_hd__buf_1 _5404_ (.A(\tree_instances[20].u_tree.read_enable ),
    .X(_2502_));
 sky130_fd_sc_hd__or2_2 _5405_ (.A(\tree_instances[20].u_tree.u_tree_weight_rom.cache_valid ),
    .B(_2502_),
    .X(_2503_));
 sky130_fd_sc_hd__buf_1 _5406_ (.A(_2503_),
    .X(_0456_));
 sky130_fd_sc_hd__inv_2 _5407_ (.A(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .Y(_2504_));
 sky130_fd_sc_hd__or2_2 _5408_ (.A(_0867_),
    .B(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .X(_2505_));
 sky130_fd_sc_hd__nand2_2 _5409_ (.A(_1488_),
    .B(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .Y(_2506_));
 sky130_fd_sc_hd__or2_2 _5410_ (.A(_0877_),
    .B(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .X(_2507_));
 sky130_fd_sc_hd__nand2_2 _5411_ (.A(_0878_),
    .B(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .Y(_2508_));
 sky130_fd_sc_hd__o21ai_2 _5412_ (.A1(_1481_),
    .A2(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .B1(\tree_instances[1].u_tree.u_tree_weight_rom.cache_valid ),
    .Y(_2509_));
 sky130_fd_sc_hd__a221o_2 _5413_ (.A1(_2505_),
    .A2(_2506_),
    .B1(_2507_),
    .B2(_2508_),
    .C1(_2509_),
    .X(_2510_));
 sky130_fd_sc_hd__o22ai_2 _5414_ (.A1(_1482_),
    .A2(_2504_),
    .B1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .B2(_1460_),
    .Y(_2511_));
 sky130_fd_sc_hd__a22o_2 _5415_ (.A1(_1461_),
    .A2(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .B2(_1459_),
    .X(_2512_));
 sky130_fd_sc_hd__a22o_2 _5416_ (.A1(_1471_),
    .A2(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .B1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .B2(_1465_),
    .X(_2513_));
 sky130_fd_sc_hd__xnor2_2 _5417_ (.A(_0868_),
    .B(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .Y(_2514_));
 sky130_fd_sc_hd__o221a_2 _5418_ (.A1(_1465_),
    .A2(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .B1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B2(_1461_),
    .C1(_2514_),
    .X(_2515_));
 sky130_fd_sc_hd__or3b_2 _5419_ (.A(_2512_),
    .B(_2513_),
    .C_N(_2515_),
    .X(_2516_));
 sky130_fd_sc_hd__a2111o_2 _5420_ (.A1(_1496_),
    .A2(_2504_),
    .B1(_2510_),
    .C1(_2511_),
    .D1(_2516_),
    .X(_2517_));
 sky130_fd_sc_hd__nand2_2 _5421_ (.A(\tree_instances[1].u_tree.read_enable ),
    .B(_2517_),
    .Y(_2518_));
 sky130_fd_sc_hd__buf_1 _5422_ (.A(_2518_),
    .X(_2519_));
 sky130_fd_sc_hd__mux2_2 _5423_ (.A0(_1496_),
    .A1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .S(_2519_),
    .X(_2520_));
 sky130_fd_sc_hd__buf_1 _5424_ (.A(_2520_),
    .X(_0457_));
 sky130_fd_sc_hd__mux2_2 _5425_ (.A0(_1492_),
    .A1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .S(_2519_),
    .X(_2521_));
 sky130_fd_sc_hd__buf_1 _5426_ (.A(_2521_),
    .X(_0458_));
 sky130_fd_sc_hd__mux2_2 _5427_ (.A0(_1494_),
    .A1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .S(_2519_),
    .X(_2522_));
 sky130_fd_sc_hd__buf_1 _5428_ (.A(_2522_),
    .X(_0459_));
 sky130_fd_sc_hd__mux2_2 _5429_ (.A0(_1497_),
    .A1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .S(_2519_),
    .X(_2523_));
 sky130_fd_sc_hd__buf_1 _5430_ (.A(_2523_),
    .X(_0460_));
 sky130_fd_sc_hd__mux2_2 _5431_ (.A0(_1495_),
    .A1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .S(_2519_),
    .X(_2524_));
 sky130_fd_sc_hd__buf_1 _5432_ (.A(_2524_),
    .X(_0461_));
 sky130_fd_sc_hd__mux2_2 _5433_ (.A0(_1480_),
    .A1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .S(_2518_),
    .X(_2525_));
 sky130_fd_sc_hd__buf_1 _5434_ (.A(_2525_),
    .X(_0462_));
 sky130_fd_sc_hd__mux2_2 _5435_ (.A0(_1489_),
    .A1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .S(_2518_),
    .X(_2526_));
 sky130_fd_sc_hd__buf_1 _5436_ (.A(_2526_),
    .X(_0463_));
 sky130_fd_sc_hd__mux2_2 _5437_ (.A0(_1498_),
    .A1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .S(_2518_),
    .X(_2527_));
 sky130_fd_sc_hd__buf_1 _5438_ (.A(_2527_),
    .X(_0464_));
 sky130_fd_sc_hd__buf_1 _5439_ (.A(_2518_),
    .X(_2528_));
 sky130_fd_sc_hd__buf_1 _5440_ (.A(_2528_),
    .X(_2529_));
 sky130_fd_sc_hd__buf_1 _5441_ (.A(\tree_instances[1].u_tree.read_enable ),
    .X(_2530_));
 sky130_fd_sc_hd__buf_1 _5442_ (.A(_2517_),
    .X(_2531_));
 sky130_fd_sc_hd__and3_2 _5443_ (.A(_2530_),
    .B(\tree_instances[1].u_tree.u_tree_weight_rom.gen_tree_1.u_tree_rom.node_data[12] ),
    .C(_2531_),
    .X(_2532_));
 sky130_fd_sc_hd__a21o_2 _5444_ (.A1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_data[12] ),
    .A2(_2529_),
    .B1(_2532_),
    .X(_0465_));
 sky130_fd_sc_hd__or3_2 _5445_ (.A(\tree_instances[1].u_tree.tree_state[1] ),
    .B(_0865_),
    .C(_1820_),
    .X(_2533_));
 sky130_fd_sc_hd__buf_1 _5446_ (.A(_2533_),
    .X(_2534_));
 sky130_fd_sc_hd__and2_2 _5447_ (.A(_1496_),
    .B(_2534_),
    .X(_2535_));
 sky130_fd_sc_hd__buf_1 _5448_ (.A(_2535_),
    .X(_0466_));
 sky130_fd_sc_hd__and2_2 _5449_ (.A(_1492_),
    .B(_2534_),
    .X(_2536_));
 sky130_fd_sc_hd__buf_1 _5450_ (.A(_2536_),
    .X(_0467_));
 sky130_fd_sc_hd__and2_2 _5451_ (.A(_1494_),
    .B(_2534_),
    .X(_2537_));
 sky130_fd_sc_hd__buf_1 _5452_ (.A(_2537_),
    .X(_0468_));
 sky130_fd_sc_hd__and2_2 _5453_ (.A(_1497_),
    .B(_2534_),
    .X(_2538_));
 sky130_fd_sc_hd__buf_1 _5454_ (.A(_2538_),
    .X(_0469_));
 sky130_fd_sc_hd__and2_2 _5455_ (.A(_1495_),
    .B(_2534_),
    .X(_2539_));
 sky130_fd_sc_hd__buf_1 _5456_ (.A(_2539_),
    .X(_0470_));
 sky130_fd_sc_hd__and2_2 _5457_ (.A(_1480_),
    .B(_2534_),
    .X(_2540_));
 sky130_fd_sc_hd__buf_1 _5458_ (.A(_2540_),
    .X(_0471_));
 sky130_fd_sc_hd__and2_2 _5459_ (.A(_1489_),
    .B(_2534_),
    .X(_2541_));
 sky130_fd_sc_hd__buf_1 _5460_ (.A(_2541_),
    .X(_0472_));
 sky130_fd_sc_hd__and2_2 _5461_ (.A(_1498_),
    .B(_2533_),
    .X(_2542_));
 sky130_fd_sc_hd__buf_1 _5462_ (.A(_2542_),
    .X(_0473_));
 sky130_fd_sc_hd__mux2_2 _5463_ (.A0(\tree_instances[20].u_tree.pipeline_frame_id[0][0] ),
    .A1(_2122_),
    .S(_0028_),
    .X(_2543_));
 sky130_fd_sc_hd__buf_1 _5464_ (.A(_2543_),
    .X(_0474_));
 sky130_fd_sc_hd__mux2_2 _5465_ (.A0(\tree_instances[20].u_tree.pipeline_frame_id[0][1] ),
    .A1(_2246_),
    .S(_0028_),
    .X(_2544_));
 sky130_fd_sc_hd__buf_1 _5466_ (.A(_2544_),
    .X(_0475_));
 sky130_fd_sc_hd__mux2_2 _5467_ (.A0(\tree_instances[20].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2125_),
    .S(_0028_),
    .X(_2545_));
 sky130_fd_sc_hd__buf_1 _5468_ (.A(_2545_),
    .X(_0476_));
 sky130_fd_sc_hd__mux2_2 _5469_ (.A0(\tree_instances[20].u_tree.pipeline_frame_id[0][3] ),
    .A1(_2249_),
    .S(_0028_),
    .X(_2546_));
 sky130_fd_sc_hd__buf_1 _5470_ (.A(_2546_),
    .X(_0477_));
 sky130_fd_sc_hd__mux2_2 _5471_ (.A0(\tree_instances[20].u_tree.pipeline_frame_id[0][4] ),
    .A1(_2251_),
    .S(_0028_),
    .X(_2547_));
 sky130_fd_sc_hd__buf_1 _5472_ (.A(_2547_),
    .X(_0478_));
 sky130_fd_sc_hd__mux2_2 _5473_ (.A0(\tree_instances[1].u_tree.current_node_data[12] ),
    .A1(\tree_instances[1].u_tree.node_data[12] ),
    .S(_0866_),
    .X(_2548_));
 sky130_fd_sc_hd__buf_1 _5474_ (.A(_2548_),
    .X(_0479_));
 sky130_fd_sc_hd__buf_1 _5475_ (.A(_0865_),
    .X(_2549_));
 sky130_fd_sc_hd__inv_2 _5476_ (.A(_0028_),
    .Y(_2550_));
 sky130_fd_sc_hd__or2b_2 _5477_ (.A(\tree_instances[20].u_tree.tree_state[1] ),
    .B_N(_2499_),
    .X(_2551_));
 sky130_fd_sc_hd__or3_2 _5478_ (.A(_0756_),
    .B(\tree_instances[20].u_tree.tree_state[1] ),
    .C(_2550_),
    .X(_2552_));
 sky130_fd_sc_hd__buf_1 _5479_ (.A(_2552_),
    .X(_2553_));
 sky130_fd_sc_hd__a21bo_2 _5480_ (.A1(_2502_),
    .A2(_2551_),
    .B1_N(_2553_),
    .X(_0480_));
 sky130_fd_sc_hd__mux2_2 _5481_ (.A0(\tree_instances[20].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[20].u_tree.pipeline_frame_id[0][0] ),
    .S(_1197_),
    .X(_2554_));
 sky130_fd_sc_hd__buf_1 _5482_ (.A(_2554_),
    .X(_0481_));
 sky130_fd_sc_hd__mux2_2 _5483_ (.A0(\tree_instances[20].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[20].u_tree.pipeline_frame_id[0][1] ),
    .S(_1197_),
    .X(_2555_));
 sky130_fd_sc_hd__buf_1 _5484_ (.A(_2555_),
    .X(_0482_));
 sky130_fd_sc_hd__mux2_2 _5485_ (.A0(\tree_instances[20].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[20].u_tree.pipeline_frame_id[0][2] ),
    .S(_1197_),
    .X(_2556_));
 sky130_fd_sc_hd__buf_1 _5486_ (.A(_2556_),
    .X(_0483_));
 sky130_fd_sc_hd__mux2_2 _5487_ (.A0(\tree_instances[20].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[20].u_tree.pipeline_frame_id[0][3] ),
    .S(_1197_),
    .X(_2557_));
 sky130_fd_sc_hd__buf_1 _5488_ (.A(_2557_),
    .X(_0484_));
 sky130_fd_sc_hd__mux2_2 _5489_ (.A0(\tree_instances[20].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[20].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[20].u_tree.tree_state[3] ),
    .X(_2558_));
 sky130_fd_sc_hd__buf_1 _5490_ (.A(_2558_),
    .X(_0485_));
 sky130_fd_sc_hd__mux2_2 _5491_ (.A0(\tree_instances[20].u_tree.prediction_out ),
    .A1(\tree_instances[20].u_tree.pipeline_prediction[0][0] ),
    .S(\tree_instances[20].u_tree.tree_state[3] ),
    .X(_2559_));
 sky130_fd_sc_hd__buf_1 _5492_ (.A(_2559_),
    .X(_0486_));
 sky130_fd_sc_hd__a22o_2 _5493_ (.A1(_1197_),
    .A2(_1198_),
    .B1(_2550_),
    .B2(\tree_instances[20].u_tree.ready_for_next ),
    .X(_0487_));
 sky130_fd_sc_hd__nand2_2 _5494_ (.A(\tree_instances[16].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[16].u_tree.tree_state[0] ),
    .Y(_2560_));
 sky130_fd_sc_hd__o2bb2a_2 _5495_ (.A1_N(_1023_),
    .A2_N(_2560_),
    .B1(_0018_),
    .B2(\tree_instances[16].u_tree.pipeline_valid[0] ),
    .X(_0488_));
 sky130_fd_sc_hd__buf_1 _5496_ (.A(\tree_instances[4].u_tree.pipeline_current_node[0][8] ),
    .X(_2561_));
 sky130_fd_sc_hd__buf_1 _5497_ (.A(_0725_),
    .X(_2562_));
 sky130_fd_sc_hd__buf_1 _5498_ (.A(_2562_),
    .X(_2563_));
 sky130_fd_sc_hd__buf_1 _5499_ (.A(_1894_),
    .X(_2564_));
 sky130_fd_sc_hd__buf_1 _5500_ (.A(_2564_),
    .X(_2565_));
 sky130_fd_sc_hd__buf_1 _5501_ (.A(_0714_),
    .X(_2566_));
 sky130_fd_sc_hd__buf_1 _5502_ (.A(_2566_),
    .X(_2567_));
 sky130_fd_sc_hd__and3_2 _5503_ (.A(_2478_),
    .B(_2484_),
    .C(_2493_),
    .X(_2568_));
 sky130_fd_sc_hd__buf_1 _5504_ (.A(_2568_),
    .X(_0490_));
 sky130_fd_sc_hd__nor2_2 _5505_ (.A(\tree_instances[11].u_tree.tree_state[3] ),
    .B(_1816_),
    .Y(_2569_));
 sky130_fd_sc_hd__o22a_2 _5506_ (.A1(\tree_instances[11].u_tree.tree_state[0] ),
    .A2(_0951_),
    .B1(_2569_),
    .B2(\tree_instances[11].u_tree.pipeline_valid[0] ),
    .X(_0491_));
 sky130_fd_sc_hd__o2bb2a_2 _5507_ (.A1_N(_0799_),
    .A2_N(_0800_),
    .B1(_0032_),
    .B2(\tree_instances[3].u_tree.pipeline_valid[0] ),
    .X(_0492_));
 sky130_fd_sc_hd__nand2_2 _5508_ (.A(\tree_instances[2].u_tree.tree_state[0] ),
    .B(_0754_),
    .Y(_2570_));
 sky130_fd_sc_hd__o2bb2a_2 _5509_ (.A1_N(_0755_),
    .A2_N(_2570_),
    .B1(_0030_),
    .B2(\tree_instances[2].u_tree.pipeline_valid[0] ),
    .X(_0493_));
 sky130_fd_sc_hd__inv_2 _5510_ (.A(\attack_votes[3] ),
    .Y(_2571_));
 sky130_fd_sc_hd__a21oi_2 _5511_ (.A1(\attack_votes[0] ),
    .A2(\attack_votes[1] ),
    .B1(\attack_votes[2] ),
    .Y(_2572_));
 sky130_fd_sc_hd__inv_2 _5512_ (.A(\attack_votes[4] ),
    .Y(_2573_));
 sky130_fd_sc_hd__o211a_2 _5513_ (.A1(_2571_),
    .A2(_2572_),
    .B1(_0000_),
    .C1(_2573_),
    .X(_2574_));
 sky130_fd_sc_hd__o21ba_2 _5514_ (.A1(prediction_out),
    .A2(_0000_),
    .B1_N(_2574_),
    .X(_0494_));
 sky130_fd_sc_hd__inv_2 _5515_ (.A(\current_voting_frame[0] ),
    .Y(_2575_));
 sky130_fd_sc_hd__buf_1 _5516_ (.A(_2575_),
    .X(_2576_));
 sky130_fd_sc_hd__nor2_2 _5517_ (.A(_2576_),
    .B(_1019_),
    .Y(_2577_));
 sky130_fd_sc_hd__a21o_2 _5518_ (.A1(frame_id_out[0]),
    .A2(_1020_),
    .B1(_2577_),
    .X(_0495_));
 sky130_fd_sc_hd__buf_1 _5519_ (.A(\current_voting_frame[1] ),
    .X(_2578_));
 sky130_fd_sc_hd__buf_1 _5520_ (.A(_2578_),
    .X(_2579_));
 sky130_fd_sc_hd__buf_1 _5521_ (.A(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__mux2_2 _5522_ (.A0(_2580_),
    .A1(frame_id_out[1]),
    .S(_1020_),
    .X(_2581_));
 sky130_fd_sc_hd__buf_1 _5523_ (.A(_2581_),
    .X(_0496_));
 sky130_fd_sc_hd__buf_1 _5524_ (.A(\current_voting_frame[2] ),
    .X(_2582_));
 sky130_fd_sc_hd__buf_1 _5525_ (.A(_2582_),
    .X(_2583_));
 sky130_fd_sc_hd__mux2_2 _5526_ (.A0(_2583_),
    .A1(frame_id_out[2]),
    .S(_1020_),
    .X(_2584_));
 sky130_fd_sc_hd__buf_1 _5527_ (.A(_2584_),
    .X(_0497_));
 sky130_fd_sc_hd__buf_1 _5528_ (.A(\current_voting_frame[3] ),
    .X(_2585_));
 sky130_fd_sc_hd__buf_1 _5529_ (.A(_2585_),
    .X(_2586_));
 sky130_fd_sc_hd__mux2_2 _5530_ (.A0(_2586_),
    .A1(frame_id_out[3]),
    .S(_1020_),
    .X(_2587_));
 sky130_fd_sc_hd__buf_1 _5531_ (.A(_2587_),
    .X(_0498_));
 sky130_fd_sc_hd__buf_1 _5532_ (.A(\current_voting_frame[4] ),
    .X(_2588_));
 sky130_fd_sc_hd__buf_1 _5533_ (.A(_2588_),
    .X(_2589_));
 sky130_fd_sc_hd__mux2_2 _5534_ (.A0(_2589_),
    .A1(frame_id_out[4]),
    .S(_1020_),
    .X(_2590_));
 sky130_fd_sc_hd__buf_1 _5535_ (.A(_2590_),
    .X(_0499_));
 sky130_fd_sc_hd__nor2_2 _5536_ (.A(\state[1] ),
    .B(_2441_),
    .Y(_2591_));
 sky130_fd_sc_hd__xor2_2 _5537_ (.A(_1827_),
    .B(_2591_),
    .X(_0500_));
 sky130_fd_sc_hd__a21oi_2 _5538_ (.A1(_1827_),
    .A2(_2591_),
    .B1(_1830_),
    .Y(_2592_));
 sky130_fd_sc_hd__and3_2 _5539_ (.A(\tree_instances[0].u_tree.frame_id_in[0] ),
    .B(\tree_instances[0].u_tree.frame_id_in[1] ),
    .C(_2591_),
    .X(_2593_));
 sky130_fd_sc_hd__nor2_2 _5540_ (.A(_2592_),
    .B(_2593_),
    .Y(_0501_));
 sky130_fd_sc_hd__xor2_2 _5541_ (.A(_1832_),
    .B(_2593_),
    .X(_0502_));
 sky130_fd_sc_hd__a21oi_2 _5542_ (.A1(_1832_),
    .A2(_2593_),
    .B1(_1835_),
    .Y(_2594_));
 sky130_fd_sc_hd__buf_1 _5543_ (.A(\tree_instances[0].u_tree.frame_id_in[2] ),
    .X(_2595_));
 sky130_fd_sc_hd__and3_2 _5544_ (.A(_2595_),
    .B(_1834_),
    .C(_2593_),
    .X(_2596_));
 sky130_fd_sc_hd__nor2_2 _5545_ (.A(_2594_),
    .B(_2596_),
    .Y(_0503_));
 sky130_fd_sc_hd__xor2_2 _5546_ (.A(_1837_),
    .B(_2596_),
    .X(_0504_));
 sky130_fd_sc_hd__nand2_2 _5547_ (.A(\attack_votes[0] ),
    .B(_1020_),
    .Y(_2597_));
 sky130_fd_sc_hd__buf_1 _5548_ (.A(_2575_),
    .X(_2598_));
 sky130_fd_sc_hd__inv_2 _5549_ (.A(_2582_),
    .Y(_2599_));
 sky130_fd_sc_hd__buf_1 _5550_ (.A(_2599_),
    .X(_2600_));
 sky130_fd_sc_hd__o2bb2a_2 _5551_ (.A1_N(_2598_),
    .A2_N(\tree_instances[20].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[20].u_tree.frame_id_out[2] ),
    .B2(_2600_),
    .X(_2601_));
 sky130_fd_sc_hd__inv_2 _5552_ (.A(\current_voting_frame[1] ),
    .Y(_2602_));
 sky130_fd_sc_hd__buf_1 _5553_ (.A(_2602_),
    .X(_2603_));
 sky130_fd_sc_hd__o2bb2a_2 _5554_ (.A1_N(_2600_),
    .A2_N(\tree_instances[20].u_tree.frame_id_out[2] ),
    .B1(\tree_instances[20].u_tree.frame_id_out[1] ),
    .B2(_2603_),
    .X(_2604_));
 sky130_fd_sc_hd__inv_2 _5555_ (.A(\current_voting_frame[3] ),
    .Y(_2605_));
 sky130_fd_sc_hd__buf_1 _5556_ (.A(_2605_),
    .X(_2606_));
 sky130_fd_sc_hd__o22a_2 _5557_ (.A1(_2598_),
    .A2(\tree_instances[20].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[20].u_tree.frame_id_out[3] ),
    .B2(_2606_),
    .X(_2607_));
 sky130_fd_sc_hd__inv_2 _5558_ (.A(\tree_instances[20].u_tree.frame_id_out[3] ),
    .Y(_2608_));
 sky130_fd_sc_hd__or2b_2 _5559_ (.A(_2578_),
    .B_N(\tree_instances[20].u_tree.frame_id_out[1] ),
    .X(_2609_));
 sky130_fd_sc_hd__buf_1 _5560_ (.A(\current_voting_frame[4] ),
    .X(_2610_));
 sky130_fd_sc_hd__xnor2_2 _5561_ (.A(_2610_),
    .B(\tree_instances[20].u_tree.frame_id_out[4] ),
    .Y(_2611_));
 sky130_fd_sc_hd__o2111a_2 _5562_ (.A1(_2585_),
    .A2(_2608_),
    .B1(_2609_),
    .C1(_2611_),
    .D1(\tree_instances[20].u_tree.prediction_valid ),
    .X(_2612_));
 sky130_fd_sc_hd__and4_2 _5563_ (.A(_2601_),
    .B(_2604_),
    .C(_2607_),
    .D(_2612_),
    .X(_2613_));
 sky130_fd_sc_hd__and2_2 _5564_ (.A(\tree_instances[20].u_tree.prediction_out ),
    .B(_2613_),
    .X(_2614_));
 sky130_fd_sc_hd__xnor2_2 _5565_ (.A(_2588_),
    .B(\tree_instances[5].u_tree.frame_id_out[4] ),
    .Y(_2615_));
 sky130_fd_sc_hd__and2_2 _5566_ (.A(_2578_),
    .B(\tree_instances[5].u_tree.frame_id_out[1] ),
    .X(_2616_));
 sky130_fd_sc_hd__nor2_2 _5567_ (.A(_2579_),
    .B(\tree_instances[5].u_tree.frame_id_out[1] ),
    .Y(_2617_));
 sky130_fd_sc_hd__o221a_2 _5568_ (.A1(_2600_),
    .A2(\tree_instances[5].u_tree.frame_id_out[2] ),
    .B1(_2616_),
    .B2(_2617_),
    .C1(\tree_instances[5].u_tree.prediction_valid ),
    .X(_2618_));
 sky130_fd_sc_hd__buf_1 _5569_ (.A(_2599_),
    .X(_2619_));
 sky130_fd_sc_hd__xor2_2 _5570_ (.A(_2585_),
    .B(\tree_instances[5].u_tree.frame_id_out[3] ),
    .X(_2620_));
 sky130_fd_sc_hd__a21oi_2 _5571_ (.A1(_2619_),
    .A2(\tree_instances[5].u_tree.frame_id_out[2] ),
    .B1(_2620_),
    .Y(_2621_));
 sky130_fd_sc_hd__buf_1 _5572_ (.A(\current_voting_frame[0] ),
    .X(_2622_));
 sky130_fd_sc_hd__xnor2_2 _5573_ (.A(_2622_),
    .B(\tree_instances[5].u_tree.frame_id_out[0] ),
    .Y(_2623_));
 sky130_fd_sc_hd__and4_2 _5574_ (.A(_2615_),
    .B(_2618_),
    .C(_2621_),
    .D(_2623_),
    .X(_2624_));
 sky130_fd_sc_hd__inv_2 _5575_ (.A(\tree_instances[3].u_tree.frame_id_out[4] ),
    .Y(_2625_));
 sky130_fd_sc_hd__xnor2_2 _5576_ (.A(_2586_),
    .B(\tree_instances[3].u_tree.frame_id_out[3] ),
    .Y(_2626_));
 sky130_fd_sc_hd__buf_1 _5577_ (.A(_2622_),
    .X(_2627_));
 sky130_fd_sc_hd__inv_2 _5578_ (.A(\tree_instances[3].u_tree.frame_id_out[0] ),
    .Y(_2628_));
 sky130_fd_sc_hd__o22a_2 _5579_ (.A1(_2575_),
    .A2(\tree_instances[3].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[3].u_tree.frame_id_out[1] ),
    .B2(_2602_),
    .X(_2629_));
 sky130_fd_sc_hd__inv_2 _5580_ (.A(\tree_instances[3].u_tree.frame_id_out[1] ),
    .Y(_2630_));
 sky130_fd_sc_hd__inv_2 _5581_ (.A(\current_voting_frame[4] ),
    .Y(_2631_));
 sky130_fd_sc_hd__xnor2_2 _5582_ (.A(_2582_),
    .B(\tree_instances[3].u_tree.frame_id_out[2] ),
    .Y(_2632_));
 sky130_fd_sc_hd__o221a_2 _5583_ (.A1(_2579_),
    .A2(_2630_),
    .B1(\tree_instances[3].u_tree.frame_id_out[4] ),
    .B2(_2631_),
    .C1(_2632_),
    .X(_2633_));
 sky130_fd_sc_hd__o211a_2 _5584_ (.A1(_2627_),
    .A2(_2628_),
    .B1(_2629_),
    .C1(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__o2111a_2 _5585_ (.A1(_2589_),
    .A2(_2625_),
    .B1(\tree_instances[3].u_tree.prediction_valid ),
    .C1(_2626_),
    .D1(_2634_),
    .X(_2635_));
 sky130_fd_sc_hd__a22o_2 _5586_ (.A1(\tree_instances[5].u_tree.prediction_out ),
    .A2(_2624_),
    .B1(_2635_),
    .B2(\tree_instances[3].u_tree.prediction_out ),
    .X(_2636_));
 sky130_fd_sc_hd__xor2_2 _5587_ (.A(_2585_),
    .B(\tree_instances[13].u_tree.frame_id_out[3] ),
    .X(_2637_));
 sky130_fd_sc_hd__a221o_2 _5588_ (.A1(_2602_),
    .A2(\tree_instances[13].u_tree.frame_id_out[1] ),
    .B1(\tree_instances[13].u_tree.frame_id_out[2] ),
    .B2(_2599_),
    .C1(_2637_),
    .X(_2638_));
 sky130_fd_sc_hd__or2b_2 _5589_ (.A(\tree_instances[13].u_tree.frame_id_out[0] ),
    .B_N(\current_voting_frame[0] ),
    .X(_2639_));
 sky130_fd_sc_hd__or2b_2 _5590_ (.A(\current_voting_frame[0] ),
    .B_N(\tree_instances[13].u_tree.frame_id_out[0] ),
    .X(_2640_));
 sky130_fd_sc_hd__o211a_2 _5591_ (.A1(_2602_),
    .A2(\tree_instances[13].u_tree.frame_id_out[1] ),
    .B1(_2639_),
    .C1(_2640_),
    .X(_2641_));
 sky130_fd_sc_hd__and2_2 _5592_ (.A(\current_voting_frame[4] ),
    .B(\tree_instances[13].u_tree.frame_id_out[4] ),
    .X(_2642_));
 sky130_fd_sc_hd__nor2_2 _5593_ (.A(_2610_),
    .B(\tree_instances[13].u_tree.frame_id_out[4] ),
    .Y(_2643_));
 sky130_fd_sc_hd__o221a_2 _5594_ (.A1(_2599_),
    .A2(\tree_instances[13].u_tree.frame_id_out[2] ),
    .B1(_2642_),
    .B2(_2643_),
    .C1(\tree_instances[13].u_tree.prediction_valid ),
    .X(_2644_));
 sky130_fd_sc_hd__and3b_2 _5595_ (.A_N(_2638_),
    .B(_2641_),
    .C(_2644_),
    .X(_2645_));
 sky130_fd_sc_hd__xnor2_2 _5596_ (.A(_2583_),
    .B(\tree_instances[1].u_tree.frame_id_out[2] ),
    .Y(_2646_));
 sky130_fd_sc_hd__xor2_2 _5597_ (.A(_2578_),
    .B(\tree_instances[1].u_tree.frame_id_out[1] ),
    .X(_2647_));
 sky130_fd_sc_hd__a221oi_2 _5598_ (.A1(_2598_),
    .A2(\tree_instances[1].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[1].u_tree.frame_id_out[3] ),
    .B2(_2606_),
    .C1(_2647_),
    .Y(_2648_));
 sky130_fd_sc_hd__or2b_2 _5599_ (.A(\tree_instances[1].u_tree.frame_id_out[3] ),
    .B_N(_2585_),
    .X(_2649_));
 sky130_fd_sc_hd__xnor2_2 _5600_ (.A(_2610_),
    .B(\tree_instances[1].u_tree.frame_id_out[4] ),
    .Y(_2650_));
 sky130_fd_sc_hd__o2111a_2 _5601_ (.A1(_2575_),
    .A2(\tree_instances[1].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[1].u_tree.prediction_valid ),
    .C1(_2649_),
    .D1(_2650_),
    .X(_2651_));
 sky130_fd_sc_hd__and3_2 _5602_ (.A(_2646_),
    .B(_2648_),
    .C(_2651_),
    .X(_2652_));
 sky130_fd_sc_hd__a22o_2 _5603_ (.A1(\tree_instances[13].u_tree.prediction_out ),
    .A2(_2645_),
    .B1(_2652_),
    .B2(\tree_instances[1].u_tree.prediction_out ),
    .X(_2653_));
 sky130_fd_sc_hd__o22a_2 _5604_ (.A1(_2576_),
    .A2(\tree_instances[8].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[8].u_tree.frame_id_out[2] ),
    .B2(_2619_),
    .X(_2654_));
 sky130_fd_sc_hd__a22o_2 _5605_ (.A1(_2575_),
    .A2(\tree_instances[8].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[8].u_tree.frame_id_out[3] ),
    .B2(_2605_),
    .X(_2655_));
 sky130_fd_sc_hd__inv_2 _5606_ (.A(\tree_instances[8].u_tree.frame_id_out[4] ),
    .Y(_2656_));
 sky130_fd_sc_hd__xor2_2 _5607_ (.A(_2578_),
    .B(\tree_instances[8].u_tree.frame_id_out[1] ),
    .X(_2657_));
 sky130_fd_sc_hd__a221o_2 _5608_ (.A1(_2600_),
    .A2(\tree_instances[8].u_tree.frame_id_out[2] ),
    .B1(_2656_),
    .B2(_2588_),
    .C1(_2657_),
    .X(_2658_));
 sky130_fd_sc_hd__buf_1 _5609_ (.A(_2605_),
    .X(_2659_));
 sky130_fd_sc_hd__o21ai_2 _5610_ (.A1(_2659_),
    .A2(\tree_instances[8].u_tree.frame_id_out[3] ),
    .B1(\tree_instances[8].u_tree.prediction_valid ),
    .Y(_2660_));
 sky130_fd_sc_hd__a2111oi_2 _5611_ (.A1(_2631_),
    .A2(\tree_instances[8].u_tree.frame_id_out[4] ),
    .B1(_2655_),
    .C1(_2658_),
    .D1(_2660_),
    .Y(_2661_));
 sky130_fd_sc_hd__and2_2 _5612_ (.A(_2610_),
    .B(\tree_instances[12].u_tree.frame_id_out[4] ),
    .X(_2662_));
 sky130_fd_sc_hd__nor2_2 _5613_ (.A(_2610_),
    .B(\tree_instances[12].u_tree.frame_id_out[4] ),
    .Y(_2663_));
 sky130_fd_sc_hd__o221a_2 _5614_ (.A1(_2600_),
    .A2(\tree_instances[12].u_tree.frame_id_out[2] ),
    .B1(_2662_),
    .B2(_2663_),
    .C1(\tree_instances[12].u_tree.prediction_valid ),
    .X(_2664_));
 sky130_fd_sc_hd__and2b_2 _5615_ (.A_N(_2585_),
    .B(\tree_instances[12].u_tree.frame_id_out[3] ),
    .X(_2665_));
 sky130_fd_sc_hd__and2b_2 _5616_ (.A_N(\tree_instances[12].u_tree.frame_id_out[3] ),
    .B(_2585_),
    .X(_2666_));
 sky130_fd_sc_hd__a211oi_2 _5617_ (.A1(_2603_),
    .A2(\tree_instances[12].u_tree.frame_id_out[1] ),
    .B1(_2665_),
    .C1(_2666_),
    .Y(_2667_));
 sky130_fd_sc_hd__inv_2 _5618_ (.A(\tree_instances[12].u_tree.frame_id_out[2] ),
    .Y(_2668_));
 sky130_fd_sc_hd__xnor2_2 _5619_ (.A(\current_voting_frame[0] ),
    .B(\tree_instances[12].u_tree.frame_id_out[0] ),
    .Y(_2669_));
 sky130_fd_sc_hd__o221a_2 _5620_ (.A1(_2602_),
    .A2(\tree_instances[12].u_tree.frame_id_out[1] ),
    .B1(_2668_),
    .B2(_2582_),
    .C1(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__and3_2 _5621_ (.A(_2664_),
    .B(_2667_),
    .C(_2670_),
    .X(_2671_));
 sky130_fd_sc_hd__a32o_2 _5622_ (.A1(\tree_instances[8].u_tree.prediction_out ),
    .A2(_2654_),
    .A3(_2661_),
    .B1(_2671_),
    .B2(\tree_instances[12].u_tree.prediction_out ),
    .X(_2672_));
 sky130_fd_sc_hd__xnor2_2 _5623_ (.A(_2585_),
    .B(\tree_instances[10].u_tree.frame_id_out[3] ),
    .Y(_2673_));
 sky130_fd_sc_hd__xor2_2 _5624_ (.A(_2610_),
    .B(\tree_instances[10].u_tree.frame_id_out[4] ),
    .X(_2674_));
 sky130_fd_sc_hd__a221oi_2 _5625_ (.A1(_2598_),
    .A2(\tree_instances[10].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[10].u_tree.frame_id_out[1] ),
    .B2(_2603_),
    .C1(_2674_),
    .Y(_2675_));
 sky130_fd_sc_hd__or2b_2 _5626_ (.A(\tree_instances[10].u_tree.frame_id_out[1] ),
    .B_N(_2578_),
    .X(_2676_));
 sky130_fd_sc_hd__xnor2_2 _5627_ (.A(_2582_),
    .B(\tree_instances[10].u_tree.frame_id_out[2] ),
    .Y(_2677_));
 sky130_fd_sc_hd__o2111a_2 _5628_ (.A1(_2575_),
    .A2(\tree_instances[10].u_tree.frame_id_out[0] ),
    .B1(_2676_),
    .C1(_2677_),
    .D1(\tree_instances[10].u_tree.prediction_valid ),
    .X(_2678_));
 sky130_fd_sc_hd__and3_2 _5629_ (.A(_2673_),
    .B(_2675_),
    .C(_2678_),
    .X(_2679_));
 sky130_fd_sc_hd__xnor2_2 _5630_ (.A(_2610_),
    .B(\tree_instances[16].u_tree.frame_id_out[4] ),
    .Y(_2680_));
 sky130_fd_sc_hd__xnor2_2 _5631_ (.A(_2582_),
    .B(\tree_instances[16].u_tree.frame_id_out[2] ),
    .Y(_2681_));
 sky130_fd_sc_hd__o2111a_2 _5632_ (.A1(_2606_),
    .A2(\tree_instances[16].u_tree.frame_id_out[3] ),
    .B1(_2680_),
    .C1(_2681_),
    .D1(\tree_instances[16].u_tree.prediction_valid ),
    .X(_2682_));
 sky130_fd_sc_hd__xnor2_2 _5633_ (.A(_2622_),
    .B(\tree_instances[16].u_tree.frame_id_out[0] ),
    .Y(_2683_));
 sky130_fd_sc_hd__and2b_2 _5634_ (.A_N(_2578_),
    .B(\tree_instances[16].u_tree.frame_id_out[1] ),
    .X(_2684_));
 sky130_fd_sc_hd__and2b_2 _5635_ (.A_N(\tree_instances[16].u_tree.frame_id_out[1] ),
    .B(_2579_),
    .X(_2685_));
 sky130_fd_sc_hd__a211oi_2 _5636_ (.A1(_2659_),
    .A2(\tree_instances[16].u_tree.frame_id_out[3] ),
    .B1(_2684_),
    .C1(_2685_),
    .Y(_2686_));
 sky130_fd_sc_hd__and3_2 _5637_ (.A(_2682_),
    .B(_2683_),
    .C(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__a22o_2 _5638_ (.A1(\tree_instances[10].u_tree.prediction_out ),
    .A2(_2679_),
    .B1(_2687_),
    .B2(\tree_instances[16].u_tree.prediction_out ),
    .X(_2688_));
 sky130_fd_sc_hd__nor3_2 _5639_ (.A(_2653_),
    .B(_2672_),
    .C(_2688_),
    .Y(_2689_));
 sky130_fd_sc_hd__or3b_2 _5640_ (.A(_2614_),
    .B(_2636_),
    .C_N(_2689_),
    .X(_2690_));
 sky130_fd_sc_hd__and2_2 _5641_ (.A(_1018_),
    .B(_2690_),
    .X(_2691_));
 sky130_fd_sc_hd__mux2_2 _5642_ (.A0(_2597_),
    .A1(\attack_votes[0] ),
    .S(_2691_),
    .X(_2692_));
 sky130_fd_sc_hd__inv_2 _5643_ (.A(_2692_),
    .Y(_0505_));
 sky130_fd_sc_hd__xor2_2 _5644_ (.A(\attack_votes[0] ),
    .B(\attack_votes[1] ),
    .X(_2693_));
 sky130_fd_sc_hd__inv_2 _5645_ (.A(\attack_votes[0] ),
    .Y(_2694_));
 sky130_fd_sc_hd__o21ba_2 _5646_ (.A1(_2694_),
    .A2(_2689_),
    .B1_N(_2636_),
    .X(_2695_));
 sky130_fd_sc_hd__a22o_2 _5647_ (.A1(_2690_),
    .A2(_2693_),
    .B1(_2695_),
    .B2(\attack_votes[1] ),
    .X(_2696_));
 sky130_fd_sc_hd__or2b_2 _5648_ (.A(_2693_),
    .B_N(_2614_),
    .X(_2697_));
 sky130_fd_sc_hd__and3_2 _5649_ (.A(\state[0] ),
    .B(_2447_),
    .C(\attack_votes[1] ),
    .X(_2698_));
 sky130_fd_sc_hd__a31o_2 _5650_ (.A1(_1018_),
    .A2(_2696_),
    .A3(_2697_),
    .B1(_2698_),
    .X(_0506_));
 sky130_fd_sc_hd__and3_2 _5651_ (.A(\attack_votes[0] ),
    .B(\attack_votes[1] ),
    .C(\attack_votes[2] ),
    .X(_2699_));
 sky130_fd_sc_hd__nor2_2 _5652_ (.A(_2572_),
    .B(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__mux2_2 _5653_ (.A0(\attack_votes[2] ),
    .A1(_2700_),
    .S(_2690_),
    .X(_2701_));
 sky130_fd_sc_hd__and3_2 _5654_ (.A(\state[0] ),
    .B(_2447_),
    .C(\attack_votes[2] ),
    .X(_2702_));
 sky130_fd_sc_hd__a21o_2 _5655_ (.A1(_1018_),
    .A2(_2701_),
    .B1(_2702_),
    .X(_0507_));
 sky130_fd_sc_hd__and3_2 _5656_ (.A(\attack_votes[3] ),
    .B(_2691_),
    .C(_2699_),
    .X(_2703_));
 sky130_fd_sc_hd__o2bb2a_2 _5657_ (.A1_N(_2691_),
    .A2_N(_2699_),
    .B1(_2571_),
    .B2(_0000_),
    .X(_2704_));
 sky130_fd_sc_hd__nor2_2 _5658_ (.A(_2703_),
    .B(_2704_),
    .Y(_0508_));
 sky130_fd_sc_hd__nor2_2 _5659_ (.A(_2573_),
    .B(_0000_),
    .Y(_2705_));
 sky130_fd_sc_hd__mux2_2 _5660_ (.A0(_2705_),
    .A1(_2573_),
    .S(_2703_),
    .X(_2706_));
 sky130_fd_sc_hd__buf_1 _5661_ (.A(_2706_),
    .X(_0509_));
 sky130_fd_sc_hd__inv_2 _5662_ (.A(\complete_votes[0] ),
    .Y(_2707_));
 sky130_fd_sc_hd__buf_1 _5663_ (.A(_2631_),
    .X(_2708_));
 sky130_fd_sc_hd__buf_1 _5664_ (.A(_2606_),
    .X(_2709_));
 sky130_fd_sc_hd__o22a_2 _5665_ (.A1(_2709_),
    .A2(\tree_instances[2].u_tree.frame_id_out[3] ),
    .B1(\tree_instances[2].u_tree.frame_id_out[4] ),
    .B2(_2708_),
    .X(_2710_));
 sky130_fd_sc_hd__a21boi_2 _5666_ (.A1(_2708_),
    .A2(\tree_instances[2].u_tree.frame_id_out[4] ),
    .B1_N(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__inv_2 _5667_ (.A(\tree_instances[2].u_tree.frame_id_out[1] ),
    .Y(_2712_));
 sky130_fd_sc_hd__buf_1 _5668_ (.A(_2603_),
    .X(_2713_));
 sky130_fd_sc_hd__buf_1 _5669_ (.A(_2619_),
    .X(_2714_));
 sky130_fd_sc_hd__o22a_2 _5670_ (.A1(_2713_),
    .A2(\tree_instances[2].u_tree.frame_id_out[1] ),
    .B1(\tree_instances[2].u_tree.frame_id_out[2] ),
    .B2(_2714_),
    .X(_2715_));
 sky130_fd_sc_hd__xor2_2 _5671_ (.A(_2627_),
    .B(\tree_instances[2].u_tree.frame_id_out[0] ),
    .X(_2716_));
 sky130_fd_sc_hd__a221oi_2 _5672_ (.A1(_2714_),
    .A2(\tree_instances[2].u_tree.frame_id_out[2] ),
    .B1(\tree_instances[2].u_tree.frame_id_out[3] ),
    .B2(_2709_),
    .C1(_2716_),
    .Y(_2717_));
 sky130_fd_sc_hd__o2111a_2 _5673_ (.A1(_2580_),
    .A2(_2712_),
    .B1(\tree_instances[2].u_tree.prediction_valid ),
    .C1(_2715_),
    .D1(_2717_),
    .X(_2718_));
 sky130_fd_sc_hd__inv_2 _5674_ (.A(\tree_instances[4].u_tree.frame_id_out[2] ),
    .Y(_2719_));
 sky130_fd_sc_hd__xnor2_2 _5675_ (.A(_2580_),
    .B(\tree_instances[4].u_tree.frame_id_out[1] ),
    .Y(_2720_));
 sky130_fd_sc_hd__inv_2 _5676_ (.A(\tree_instances[4].u_tree.frame_id_out[0] ),
    .Y(_2721_));
 sky130_fd_sc_hd__and2_2 _5677_ (.A(_2589_),
    .B(\tree_instances[4].u_tree.frame_id_out[4] ),
    .X(_2722_));
 sky130_fd_sc_hd__nor2_2 _5678_ (.A(_2589_),
    .B(\tree_instances[4].u_tree.frame_id_out[4] ),
    .Y(_2723_));
 sky130_fd_sc_hd__xnor2_2 _5679_ (.A(_2586_),
    .B(\tree_instances[4].u_tree.frame_id_out[3] ),
    .Y(_2724_));
 sky130_fd_sc_hd__o221a_2 _5680_ (.A1(_2576_),
    .A2(\tree_instances[4].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[4].u_tree.frame_id_out[2] ),
    .B2(_2714_),
    .C1(_2724_),
    .X(_2725_));
 sky130_fd_sc_hd__o221a_2 _5681_ (.A1(_2627_),
    .A2(_2721_),
    .B1(_2722_),
    .B2(_2723_),
    .C1(_2725_),
    .X(_2726_));
 sky130_fd_sc_hd__o2111a_2 _5682_ (.A1(_2583_),
    .A2(_2719_),
    .B1(\tree_instances[4].u_tree.prediction_valid ),
    .C1(_2720_),
    .D1(_2726_),
    .X(_2727_));
 sky130_fd_sc_hd__a211oi_2 _5683_ (.A1(_2711_),
    .A2(_2718_),
    .B1(_2635_),
    .C1(_2727_),
    .Y(_2728_));
 sky130_fd_sc_hd__inv_2 _5684_ (.A(_2728_),
    .Y(_2729_));
 sky130_fd_sc_hd__inv_2 _5685_ (.A(\tree_instances[9].u_tree.frame_id_out[1] ),
    .Y(_2730_));
 sky130_fd_sc_hd__o22a_2 _5686_ (.A1(_2713_),
    .A2(\tree_instances[9].u_tree.frame_id_out[1] ),
    .B1(\tree_instances[9].u_tree.frame_id_out[4] ),
    .B2(_2708_),
    .X(_2731_));
 sky130_fd_sc_hd__inv_2 _5687_ (.A(\tree_instances[9].u_tree.frame_id_out[0] ),
    .Y(_2732_));
 sky130_fd_sc_hd__xor2_2 _5688_ (.A(_2582_),
    .B(\tree_instances[9].u_tree.frame_id_out[2] ),
    .X(_2733_));
 sky130_fd_sc_hd__a221o_2 _5689_ (.A1(_2622_),
    .A2(_2732_),
    .B1(\tree_instances[9].u_tree.frame_id_out[4] ),
    .B2(_2631_),
    .C1(_2733_),
    .X(_2734_));
 sky130_fd_sc_hd__a22o_2 _5690_ (.A1(_2598_),
    .A2(\tree_instances[9].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[9].u_tree.frame_id_out[3] ),
    .B2(_2659_),
    .X(_2735_));
 sky130_fd_sc_hd__o21ai_2 _5691_ (.A1(_2659_),
    .A2(\tree_instances[9].u_tree.frame_id_out[3] ),
    .B1(\tree_instances[9].u_tree.prediction_valid ),
    .Y(_2736_));
 sky130_fd_sc_hd__nor3_2 _5692_ (.A(_2734_),
    .B(_2735_),
    .C(_2736_),
    .Y(_2737_));
 sky130_fd_sc_hd__o211a_2 _5693_ (.A1(_2580_),
    .A2(_2730_),
    .B1(_2731_),
    .C1(_2737_),
    .X(_2738_));
 sky130_fd_sc_hd__inv_2 _5694_ (.A(\tree_instances[17].u_tree.frame_id_out[0] ),
    .Y(_2739_));
 sky130_fd_sc_hd__o22a_2 _5695_ (.A1(_2576_),
    .A2(\tree_instances[17].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[17].u_tree.frame_id_out[1] ),
    .B2(_2713_),
    .X(_2740_));
 sky130_fd_sc_hd__xor2_2 _5696_ (.A(_2582_),
    .B(\tree_instances[17].u_tree.frame_id_out[2] ),
    .X(_2741_));
 sky130_fd_sc_hd__a221oi_2 _5697_ (.A1(_2603_),
    .A2(\tree_instances[17].u_tree.frame_id_out[1] ),
    .B1(\tree_instances[17].u_tree.frame_id_out[3] ),
    .B2(_2659_),
    .C1(_2741_),
    .Y(_2742_));
 sky130_fd_sc_hd__xnor2_2 _5698_ (.A(_2588_),
    .B(\tree_instances[17].u_tree.frame_id_out[4] ),
    .Y(_2743_));
 sky130_fd_sc_hd__o2111a_2 _5699_ (.A1(_2659_),
    .A2(\tree_instances[17].u_tree.frame_id_out[3] ),
    .B1(_2742_),
    .C1(_2743_),
    .D1(\tree_instances[17].u_tree.prediction_valid ),
    .X(_2744_));
 sky130_fd_sc_hd__o211a_2 _5700_ (.A1(_2627_),
    .A2(_2739_),
    .B1(_2740_),
    .C1(_2744_),
    .X(_2745_));
 sky130_fd_sc_hd__inv_2 _5701_ (.A(\tree_instances[0].u_tree.frame_id_out[2] ),
    .Y(_2746_));
 sky130_fd_sc_hd__xnor2_2 _5702_ (.A(\tree_instances[0].u_tree.frame_id_out[4] ),
    .B(_2588_),
    .Y(_2747_));
 sky130_fd_sc_hd__o221a_2 _5703_ (.A1(_2746_),
    .A2(_2583_),
    .B1(\tree_instances[0].u_tree.frame_id_out[3] ),
    .B2(_2659_),
    .C1(_2747_),
    .X(_2748_));
 sky130_fd_sc_hd__inv_2 _5704_ (.A(\tree_instances[0].u_tree.frame_id_out[0] ),
    .Y(_2749_));
 sky130_fd_sc_hd__o2bb2a_2 _5705_ (.A1_N(\tree_instances[0].u_tree.frame_id_out[3] ),
    .A2_N(_2606_),
    .B1(\tree_instances[0].u_tree.frame_id_out[0] ),
    .B2(_2598_),
    .X(_2750_));
 sky130_fd_sc_hd__and2_2 _5706_ (.A(\tree_instances[0].u_tree.frame_id_out[1] ),
    .B(_2578_),
    .X(_2751_));
 sky130_fd_sc_hd__nor2_2 _5707_ (.A(\tree_instances[0].u_tree.frame_id_out[1] ),
    .B(_2579_),
    .Y(_2752_));
 sky130_fd_sc_hd__o221a_2 _5708_ (.A1(\tree_instances[0].u_tree.frame_id_out[2] ),
    .A2(_2600_),
    .B1(_2751_),
    .B2(_2752_),
    .C1(\tree_instances[0].u_tree.prediction_valid ),
    .X(_2753_));
 sky130_fd_sc_hd__o211a_2 _5709_ (.A1(_2749_),
    .A2(_2627_),
    .B1(_2750_),
    .C1(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__a211o_2 _5710_ (.A1(_2748_),
    .A2(_2754_),
    .B1(_2652_),
    .C1(_2679_),
    .X(_2755_));
 sky130_fd_sc_hd__a22oi_2 _5711_ (.A1(_2713_),
    .A2(\tree_instances[18].u_tree.frame_id_out[1] ),
    .B1(\tree_instances[18].u_tree.frame_id_out[2] ),
    .B2(_2714_),
    .Y(_2756_));
 sky130_fd_sc_hd__inv_2 _5712_ (.A(\tree_instances[18].u_tree.frame_id_out[3] ),
    .Y(_2757_));
 sky130_fd_sc_hd__and2_2 _5713_ (.A(_2622_),
    .B(\tree_instances[18].u_tree.frame_id_out[0] ),
    .X(_2758_));
 sky130_fd_sc_hd__nor2_2 _5714_ (.A(_2622_),
    .B(\tree_instances[18].u_tree.frame_id_out[0] ),
    .Y(_2759_));
 sky130_fd_sc_hd__xnor2_2 _5715_ (.A(_2588_),
    .B(\tree_instances[18].u_tree.frame_id_out[4] ),
    .Y(_2760_));
 sky130_fd_sc_hd__o221a_2 _5716_ (.A1(_2606_),
    .A2(\tree_instances[18].u_tree.frame_id_out[3] ),
    .B1(_2758_),
    .B2(_2759_),
    .C1(_2760_),
    .X(_2761_));
 sky130_fd_sc_hd__o221a_2 _5717_ (.A1(_2619_),
    .A2(\tree_instances[18].u_tree.frame_id_out[2] ),
    .B1(_2757_),
    .B2(_2586_),
    .C1(_2761_),
    .X(_2762_));
 sky130_fd_sc_hd__o2111a_2 _5718_ (.A1(_2713_),
    .A2(\tree_instances[18].u_tree.frame_id_out[1] ),
    .B1(_2756_),
    .C1(_2762_),
    .D1(\tree_instances[18].u_tree.prediction_valid ),
    .X(_2763_));
 sky130_fd_sc_hd__or4_2 _5719_ (.A(_2738_),
    .B(_2745_),
    .C(_2755_),
    .D(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__a2bb2o_2 _5720_ (.A1_N(_2708_),
    .A2_N(\tree_instances[15].u_tree.frame_id_out[4] ),
    .B1(\tree_instances[15].u_tree.frame_id_out[3] ),
    .B2(_2709_),
    .X(_2765_));
 sky130_fd_sc_hd__a21o_2 _5721_ (.A1(_2708_),
    .A2(\tree_instances[15].u_tree.frame_id_out[4] ),
    .B1(_2765_),
    .X(_2766_));
 sky130_fd_sc_hd__nor2_2 _5722_ (.A(_2714_),
    .B(\tree_instances[15].u_tree.frame_id_out[2] ),
    .Y(_2767_));
 sky130_fd_sc_hd__a22o_2 _5723_ (.A1(_2576_),
    .A2(\tree_instances[15].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[15].u_tree.frame_id_out[2] ),
    .B2(_2714_),
    .X(_2768_));
 sky130_fd_sc_hd__o2bb2a_2 _5724_ (.A1_N(_2603_),
    .A2_N(\tree_instances[15].u_tree.frame_id_out[1] ),
    .B1(\tree_instances[15].u_tree.frame_id_out[0] ),
    .B2(_2598_),
    .X(_2769_));
 sky130_fd_sc_hd__o221a_2 _5725_ (.A1(_2713_),
    .A2(\tree_instances[15].u_tree.frame_id_out[1] ),
    .B1(\tree_instances[15].u_tree.frame_id_out[3] ),
    .B2(_2709_),
    .C1(_2769_),
    .X(_2770_));
 sky130_fd_sc_hd__or4bb_2 _5726_ (.A(_2767_),
    .B(_2768_),
    .C_N(\tree_instances[15].u_tree.prediction_valid ),
    .D_N(_2770_),
    .X(_2771_));
 sky130_fd_sc_hd__inv_2 _5727_ (.A(\tree_instances[19].u_tree.frame_id_out[4] ),
    .Y(_2772_));
 sky130_fd_sc_hd__a22o_2 _5728_ (.A1(_2709_),
    .A2(\tree_instances[19].u_tree.frame_id_out[3] ),
    .B1(_2772_),
    .B2(_2589_),
    .X(_2773_));
 sky130_fd_sc_hd__a21bo_2 _5729_ (.A1(_2714_),
    .A2(\tree_instances[19].u_tree.frame_id_out[2] ),
    .B1_N(\tree_instances[19].u_tree.prediction_valid ),
    .X(_2774_));
 sky130_fd_sc_hd__o22a_2 _5730_ (.A1(_2576_),
    .A2(\tree_instances[19].u_tree.frame_id_out[0] ),
    .B1(_2772_),
    .B2(_2588_),
    .X(_2775_));
 sky130_fd_sc_hd__inv_2 _5731_ (.A(\tree_instances[19].u_tree.frame_id_out[0] ),
    .Y(_2776_));
 sky130_fd_sc_hd__xnor2_2 _5732_ (.A(_2579_),
    .B(\tree_instances[19].u_tree.frame_id_out[1] ),
    .Y(_2777_));
 sky130_fd_sc_hd__o221a_2 _5733_ (.A1(_2627_),
    .A2(_2776_),
    .B1(\tree_instances[19].u_tree.frame_id_out[2] ),
    .B2(_2619_),
    .C1(_2777_),
    .X(_2778_));
 sky130_fd_sc_hd__o211a_2 _5734_ (.A1(_2709_),
    .A2(\tree_instances[19].u_tree.frame_id_out[3] ),
    .B1(_2775_),
    .C1(_2778_),
    .X(_2779_));
 sky130_fd_sc_hd__or3b_2 _5735_ (.A(_2773_),
    .B(_2774_),
    .C_N(_2779_),
    .X(_2780_));
 sky130_fd_sc_hd__o2bb2a_2 _5736_ (.A1_N(_2708_),
    .A2_N(\tree_instances[14].u_tree.frame_id_out[4] ),
    .B1(\tree_instances[14].u_tree.frame_id_out[2] ),
    .B2(_2714_),
    .X(_2781_));
 sky130_fd_sc_hd__inv_2 _5737_ (.A(\tree_instances[14].u_tree.frame_id_out[3] ),
    .Y(_2782_));
 sky130_fd_sc_hd__inv_2 _5738_ (.A(\tree_instances[14].u_tree.frame_id_out[2] ),
    .Y(_2783_));
 sky130_fd_sc_hd__xnor2_2 _5739_ (.A(_2579_),
    .B(\tree_instances[14].u_tree.frame_id_out[1] ),
    .Y(_2784_));
 sky130_fd_sc_hd__o221a_2 _5740_ (.A1(_2583_),
    .A2(_2783_),
    .B1(\tree_instances[14].u_tree.frame_id_out[4] ),
    .B2(_2708_),
    .C1(_2784_),
    .X(_2785_));
 sky130_fd_sc_hd__xnor2_2 _5741_ (.A(_2627_),
    .B(\tree_instances[14].u_tree.frame_id_out[0] ),
    .Y(_2786_));
 sky130_fd_sc_hd__o211a_2 _5742_ (.A1(_2709_),
    .A2(\tree_instances[14].u_tree.frame_id_out[3] ),
    .B1(_2786_),
    .C1(\tree_instances[14].u_tree.prediction_valid ),
    .X(_2787_));
 sky130_fd_sc_hd__o211a_2 _5743_ (.A1(_2586_),
    .A2(_2782_),
    .B1(_2785_),
    .C1(_2787_),
    .X(_2788_));
 sky130_fd_sc_hd__and2b_2 _5744_ (.A_N(\tree_instances[11].u_tree.frame_id_out[1] ),
    .B(_2579_),
    .X(_2789_));
 sky130_fd_sc_hd__and2b_2 _5745_ (.A_N(_2580_),
    .B(\tree_instances[11].u_tree.frame_id_out[1] ),
    .X(_2790_));
 sky130_fd_sc_hd__a211oi_2 _5746_ (.A1(_2576_),
    .A2(\tree_instances[11].u_tree.frame_id_out[0] ),
    .B1(_2789_),
    .C1(_2790_),
    .Y(_2791_));
 sky130_fd_sc_hd__xnor2_2 _5747_ (.A(_2586_),
    .B(\tree_instances[11].u_tree.frame_id_out[3] ),
    .Y(_2792_));
 sky130_fd_sc_hd__o221a_2 _5748_ (.A1(_2576_),
    .A2(\tree_instances[11].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[11].u_tree.frame_id_out[2] ),
    .B2(_2619_),
    .C1(_2792_),
    .X(_2793_));
 sky130_fd_sc_hd__inv_2 _5749_ (.A(\tree_instances[11].u_tree.frame_id_out[2] ),
    .Y(_2794_));
 sky130_fd_sc_hd__and2_2 _5750_ (.A(_2588_),
    .B(\tree_instances[11].u_tree.frame_id_out[4] ),
    .X(_2795_));
 sky130_fd_sc_hd__nor2_2 _5751_ (.A(_2589_),
    .B(\tree_instances[11].u_tree.frame_id_out[4] ),
    .Y(_2796_));
 sky130_fd_sc_hd__o221a_2 _5752_ (.A1(_2583_),
    .A2(_2794_),
    .B1(_2795_),
    .B2(_2796_),
    .C1(\tree_instances[11].u_tree.prediction_valid ),
    .X(_2797_));
 sky130_fd_sc_hd__and3_2 _5753_ (.A(_2791_),
    .B(_2793_),
    .C(_2797_),
    .X(_2798_));
 sky130_fd_sc_hd__a21oi_2 _5754_ (.A1(_2781_),
    .A2(_2788_),
    .B1(_2798_),
    .Y(_2799_));
 sky130_fd_sc_hd__o211ai_2 _5755_ (.A1(_2766_),
    .A2(_2771_),
    .B1(_2780_),
    .C1(_2799_),
    .Y(_2800_));
 sky130_fd_sc_hd__inv_2 _5756_ (.A(\tree_instances[6].u_tree.frame_id_out[1] ),
    .Y(_2801_));
 sky130_fd_sc_hd__and2_2 _5757_ (.A(_2622_),
    .B(\tree_instances[6].u_tree.frame_id_out[0] ),
    .X(_2802_));
 sky130_fd_sc_hd__nor2_2 _5758_ (.A(_2622_),
    .B(\tree_instances[6].u_tree.frame_id_out[0] ),
    .Y(_2803_));
 sky130_fd_sc_hd__o221a_2 _5759_ (.A1(_2580_),
    .A2(_2801_),
    .B1(_2802_),
    .B2(_2803_),
    .C1(\tree_instances[6].u_tree.prediction_valid ),
    .X(_2804_));
 sky130_fd_sc_hd__nand2_2 _5760_ (.A(_2659_),
    .B(\tree_instances[6].u_tree.frame_id_out[3] ),
    .Y(_2805_));
 sky130_fd_sc_hd__o221a_2 _5761_ (.A1(_2603_),
    .A2(\tree_instances[6].u_tree.frame_id_out[1] ),
    .B1(\tree_instances[6].u_tree.frame_id_out[4] ),
    .B2(_2708_),
    .C1(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__inv_2 _5762_ (.A(\tree_instances[6].u_tree.frame_id_out[4] ),
    .Y(_2807_));
 sky130_fd_sc_hd__o2bb2a_2 _5763_ (.A1_N(_2600_),
    .A2_N(\tree_instances[6].u_tree.frame_id_out[2] ),
    .B1(\tree_instances[6].u_tree.frame_id_out[3] ),
    .B2(_2606_),
    .X(_2808_));
 sky130_fd_sc_hd__o221a_2 _5764_ (.A1(_2619_),
    .A2(\tree_instances[6].u_tree.frame_id_out[2] ),
    .B1(_2807_),
    .B2(_2589_),
    .C1(_2808_),
    .X(_2809_));
 sky130_fd_sc_hd__and3_2 _5765_ (.A(_2804_),
    .B(_2806_),
    .C(_2809_),
    .X(_2810_));
 sky130_fd_sc_hd__a22o_2 _5766_ (.A1(_2619_),
    .A2(\tree_instances[7].u_tree.frame_id_out[2] ),
    .B1(\tree_instances[7].u_tree.frame_id_out[3] ),
    .B2(_2606_),
    .X(_2811_));
 sky130_fd_sc_hd__o21ba_2 _5767_ (.A1(_2709_),
    .A2(\tree_instances[7].u_tree.frame_id_out[3] ),
    .B1_N(_2811_),
    .X(_2812_));
 sky130_fd_sc_hd__xnor2_2 _5768_ (.A(_2610_),
    .B(\tree_instances[7].u_tree.frame_id_out[4] ),
    .Y(_2813_));
 sky130_fd_sc_hd__o221a_2 _5769_ (.A1(_2575_),
    .A2(\tree_instances[7].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[7].u_tree.frame_id_out[2] ),
    .B2(_2600_),
    .C1(_2813_),
    .X(_2814_));
 sky130_fd_sc_hd__a22oi_2 _5770_ (.A1(_2598_),
    .A2(\tree_instances[7].u_tree.frame_id_out[0] ),
    .B1(\tree_instances[7].u_tree.frame_id_out[1] ),
    .B2(_2603_),
    .Y(_2815_));
 sky130_fd_sc_hd__o2111a_2 _5771_ (.A1(_2713_),
    .A2(\tree_instances[7].u_tree.frame_id_out[1] ),
    .B1(_2814_),
    .C1(_2815_),
    .D1(\tree_instances[7].u_tree.prediction_valid ),
    .X(_2816_));
 sky130_fd_sc_hd__a211o_2 _5772_ (.A1(_2812_),
    .A2(_2816_),
    .B1(_2624_),
    .C1(_2613_),
    .X(_2817_));
 sky130_fd_sc_hd__a211o_2 _5773_ (.A1(_2654_),
    .A2(_2661_),
    .B1(_2671_),
    .C1(_2645_),
    .X(_2818_));
 sky130_fd_sc_hd__or4_2 _5774_ (.A(_2687_),
    .B(_2810_),
    .C(_2817_),
    .D(_2818_),
    .X(_2819_));
 sky130_fd_sc_hd__or3_2 _5775_ (.A(_2764_),
    .B(_2800_),
    .C(_2819_),
    .X(_2820_));
 sky130_fd_sc_hd__nor2_2 _5776_ (.A(_2729_),
    .B(_2820_),
    .Y(_2821_));
 sky130_fd_sc_hd__a2bb2o_2 _5777_ (.A1_N(_2447_),
    .A2_N(_2821_),
    .B1(_1020_),
    .B2(\complete_votes[0] ),
    .X(_2822_));
 sky130_fd_sc_hd__o31a_2 _5778_ (.A1(_2447_),
    .A2(_2707_),
    .A3(_2821_),
    .B1(_2822_),
    .X(_0510_));
 sky130_fd_sc_hd__inv_2 _5779_ (.A(\complete_votes[1] ),
    .Y(_2823_));
 sky130_fd_sc_hd__o32a_2 _5780_ (.A1(_2447_),
    .A2(_2707_),
    .A3(_2821_),
    .B1(_0000_),
    .B2(_2823_),
    .X(_2824_));
 sky130_fd_sc_hd__o2111a_2 _5781_ (.A1(_2729_),
    .A2(_2820_),
    .B1(_1018_),
    .C1(\complete_votes[1] ),
    .D1(\complete_votes[0] ),
    .X(_2825_));
 sky130_fd_sc_hd__nor2_2 _5782_ (.A(_2824_),
    .B(_2825_),
    .Y(_0511_));
 sky130_fd_sc_hd__inv_2 _5783_ (.A(\complete_votes[2] ),
    .Y(_2826_));
 sky130_fd_sc_hd__nor2_2 _5784_ (.A(_2826_),
    .B(_0000_),
    .Y(_2827_));
 sky130_fd_sc_hd__mux2_2 _5785_ (.A0(_2827_),
    .A1(_2826_),
    .S(_2825_),
    .X(_2828_));
 sky130_fd_sc_hd__buf_1 _5786_ (.A(_2828_),
    .X(_0512_));
 sky130_fd_sc_hd__nor2_2 _5787_ (.A(_2823_),
    .B(_2444_),
    .Y(_2829_));
 sky130_fd_sc_hd__xnor2_2 _5788_ (.A(\complete_votes[3] ),
    .B(_2829_),
    .Y(_2830_));
 sky130_fd_sc_hd__a2bb2o_2 _5789_ (.A1_N(_2821_),
    .A2_N(_2830_),
    .B1(\complete_votes[3] ),
    .B2(_2728_),
    .X(_2831_));
 sky130_fd_sc_hd__a21oi_2 _5790_ (.A1(_2820_),
    .A2(_2830_),
    .B1(_2447_),
    .Y(_2832_));
 sky130_fd_sc_hd__a32o_2 _5791_ (.A1(\state[0] ),
    .A2(_2447_),
    .A3(\complete_votes[3] ),
    .B1(_2831_),
    .B2(_2832_),
    .X(_0513_));
 sky130_fd_sc_hd__nor2_2 _5792_ (.A(_2443_),
    .B(_1021_),
    .Y(_2833_));
 sky130_fd_sc_hd__o2111a_2 _5793_ (.A1(_2729_),
    .A2(_2820_),
    .B1(_2829_),
    .C1(\complete_votes[3] ),
    .D1(_1018_),
    .X(_2834_));
 sky130_fd_sc_hd__mux2_2 _5794_ (.A0(_2833_),
    .A1(_2443_),
    .S(_2834_),
    .X(_2835_));
 sky130_fd_sc_hd__buf_1 _5795_ (.A(_2835_),
    .X(_0514_));
 sky130_fd_sc_hd__nor2_2 _5796_ (.A(_2627_),
    .B(_0000_),
    .Y(_2836_));
 sky130_fd_sc_hd__nor2_2 _5797_ (.A(_2577_),
    .B(_2836_),
    .Y(_0515_));
 sky130_fd_sc_hd__xnor2_2 _5798_ (.A(_2713_),
    .B(_2577_),
    .Y(_0516_));
 sky130_fd_sc_hd__and3_2 _5799_ (.A(_2580_),
    .B(_2583_),
    .C(_2577_),
    .X(_2837_));
 sky130_fd_sc_hd__a21oi_2 _5800_ (.A1(_2580_),
    .A2(_2577_),
    .B1(_2583_),
    .Y(_2838_));
 sky130_fd_sc_hd__nor2_2 _5801_ (.A(_2837_),
    .B(_2838_),
    .Y(_0517_));
 sky130_fd_sc_hd__nand2_2 _5802_ (.A(_2586_),
    .B(_2837_),
    .Y(_2839_));
 sky130_fd_sc_hd__or2_2 _5803_ (.A(_2586_),
    .B(_2837_),
    .X(_2840_));
 sky130_fd_sc_hd__and2_2 _5804_ (.A(_2839_),
    .B(_2840_),
    .X(_2841_));
 sky130_fd_sc_hd__buf_1 _5805_ (.A(_2841_),
    .X(_0518_));
 sky130_fd_sc_hd__xnor2_2 _5806_ (.A(_2589_),
    .B(_2839_),
    .Y(_0519_));
 sky130_fd_sc_hd__mux2_2 _5807_ (.A0(\tree_instances[0].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1826_),
    .S(_0004_),
    .X(_2842_));
 sky130_fd_sc_hd__buf_1 _5808_ (.A(_2842_),
    .X(_0520_));
 sky130_fd_sc_hd__mux2_2 _5809_ (.A0(\tree_instances[0].u_tree.pipeline_frame_id[0][1] ),
    .A1(_2246_),
    .S(_0004_),
    .X(_2843_));
 sky130_fd_sc_hd__buf_1 _5810_ (.A(_2843_),
    .X(_0521_));
 sky130_fd_sc_hd__mux2_2 _5811_ (.A0(\tree_instances[0].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2595_),
    .S(_0004_),
    .X(_2844_));
 sky130_fd_sc_hd__buf_1 _5812_ (.A(_2844_),
    .X(_0522_));
 sky130_fd_sc_hd__mux2_2 _5813_ (.A0(\tree_instances[0].u_tree.pipeline_frame_id[0][3] ),
    .A1(_2249_),
    .S(_0004_),
    .X(_2845_));
 sky130_fd_sc_hd__buf_1 _5814_ (.A(_2845_),
    .X(_0523_));
 sky130_fd_sc_hd__mux2_2 _5815_ (.A0(\tree_instances[0].u_tree.pipeline_frame_id[0][4] ),
    .A1(_2251_),
    .S(_0004_),
    .X(_2846_));
 sky130_fd_sc_hd__buf_1 _5816_ (.A(_2846_),
    .X(_0524_));
 sky130_fd_sc_hd__mux2_2 _5817_ (.A0(\tree_instances[0].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[0].u_tree.pipeline_frame_id[0][0] ),
    .S(_0737_),
    .X(_2847_));
 sky130_fd_sc_hd__buf_1 _5818_ (.A(_2847_),
    .X(_0525_));
 sky130_fd_sc_hd__mux2_2 _5819_ (.A0(\tree_instances[0].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[0].u_tree.pipeline_frame_id[0][1] ),
    .S(_0737_),
    .X(_2848_));
 sky130_fd_sc_hd__buf_1 _5820_ (.A(_2848_),
    .X(_0526_));
 sky130_fd_sc_hd__mux2_2 _5821_ (.A0(\tree_instances[0].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[0].u_tree.pipeline_frame_id[0][2] ),
    .S(_0737_),
    .X(_2849_));
 sky130_fd_sc_hd__buf_1 _5822_ (.A(_2849_),
    .X(_0527_));
 sky130_fd_sc_hd__mux2_2 _5823_ (.A0(\tree_instances[0].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[0].u_tree.pipeline_frame_id[0][3] ),
    .S(_0737_),
    .X(_2850_));
 sky130_fd_sc_hd__buf_1 _5824_ (.A(_2850_),
    .X(_0528_));
 sky130_fd_sc_hd__mux2_2 _5825_ (.A0(\tree_instances[0].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[0].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[0].u_tree.tree_state[3] ),
    .X(_2851_));
 sky130_fd_sc_hd__buf_1 _5826_ (.A(_2851_),
    .X(_0529_));
 sky130_fd_sc_hd__a22o_2 _5827_ (.A1(_0737_),
    .A2(_2495_),
    .B1(_1818_),
    .B2(\tree_instances[0].u_tree.ready_for_next ),
    .X(_0530_));
 sky130_fd_sc_hd__nor2_2 _5828_ (.A(_1932_),
    .B(_1968_),
    .Y(_2852_));
 sky130_fd_sc_hd__buf_1 _5829_ (.A(_2852_),
    .X(_2853_));
 sky130_fd_sc_hd__a221o_2 _5830_ (.A1(_1934_),
    .A2(\tree_instances[8].u_tree.node_data[12] ),
    .B1(_2853_),
    .B2(\tree_instances[8].u_tree.u_tree_weight_rom.cached_data[12] ),
    .C1(_1967_),
    .X(_0531_));
 sky130_fd_sc_hd__a22o_2 _5831_ (.A1(\tree_instances[1].u_tree.tree_state[1] ),
    .A2(\tree_instances[1].u_tree.current_node_data[12] ),
    .B1(\tree_instances[1].u_tree.node_data[12] ),
    .B2(_2549_),
    .X(_2854_));
 sky130_fd_sc_hd__nand2_2 _5832_ (.A(\tree_instances[1].u_tree.tree_state[0] ),
    .B(_1226_),
    .Y(_2855_));
 sky130_fd_sc_hd__or3_2 _5833_ (.A(\tree_instances[1].u_tree.tree_state[1] ),
    .B(\tree_instances[1].u_tree.tree_state[0] ),
    .C(\tree_instances[1].u_tree.tree_state[2] ),
    .X(_2856_));
 sky130_fd_sc_hd__o211a_2 _5834_ (.A1(_1821_),
    .A2(_0883_),
    .B1(_2855_),
    .C1(_2856_),
    .X(_2857_));
 sky130_fd_sc_hd__mux2_2 _5835_ (.A0(\tree_instances[1].u_tree.pipeline_prediction[0][0] ),
    .A1(_2854_),
    .S(_2857_),
    .X(_2858_));
 sky130_fd_sc_hd__buf_1 _5836_ (.A(_2858_),
    .X(_0532_));
 sky130_fd_sc_hd__a21o_2 _5837_ (.A1(_2530_),
    .A2(_2531_),
    .B1(\tree_instances[1].u_tree.u_tree_weight_rom.cache_valid ),
    .X(_0533_));
 sky130_fd_sc_hd__and2_2 _5838_ (.A(_1527_),
    .B(_2427_),
    .X(_2859_));
 sky130_fd_sc_hd__buf_1 _5839_ (.A(_2859_),
    .X(_0534_));
 sky130_fd_sc_hd__and2_2 _5840_ (.A(_1512_),
    .B(_2427_),
    .X(_2860_));
 sky130_fd_sc_hd__buf_1 _5841_ (.A(_2860_),
    .X(_0535_));
 sky130_fd_sc_hd__and2_2 _5842_ (.A(_1516_),
    .B(_2427_),
    .X(_2861_));
 sky130_fd_sc_hd__buf_1 _5843_ (.A(_2861_),
    .X(_0536_));
 sky130_fd_sc_hd__and2_2 _5844_ (.A(_1519_),
    .B(_2427_),
    .X(_2862_));
 sky130_fd_sc_hd__buf_1 _5845_ (.A(_2862_),
    .X(_0537_));
 sky130_fd_sc_hd__and2_2 _5846_ (.A(_1526_),
    .B(_2427_),
    .X(_2863_));
 sky130_fd_sc_hd__buf_1 _5847_ (.A(_2863_),
    .X(_0538_));
 sky130_fd_sc_hd__and2_2 _5848_ (.A(_1525_),
    .B(_2427_),
    .X(_2864_));
 sky130_fd_sc_hd__buf_1 _5849_ (.A(_2864_),
    .X(_0539_));
 sky130_fd_sc_hd__and2_2 _5850_ (.A(_1510_),
    .B(_2427_),
    .X(_2865_));
 sky130_fd_sc_hd__buf_1 _5851_ (.A(_2865_),
    .X(_0540_));
 sky130_fd_sc_hd__and2_2 _5852_ (.A(_1522_),
    .B(_2426_),
    .X(_2866_));
 sky130_fd_sc_hd__buf_1 _5853_ (.A(_2866_),
    .X(_0541_));
 sky130_fd_sc_hd__mux2_2 _5854_ (.A0(\tree_instances[1].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1826_),
    .S(_0026_),
    .X(_2867_));
 sky130_fd_sc_hd__buf_1 _5855_ (.A(_2867_),
    .X(_0542_));
 sky130_fd_sc_hd__mux2_2 _5856_ (.A0(\tree_instances[1].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1829_),
    .S(_0026_),
    .X(_2868_));
 sky130_fd_sc_hd__buf_1 _5857_ (.A(_2868_),
    .X(_0543_));
 sky130_fd_sc_hd__mux2_2 _5858_ (.A0(\tree_instances[1].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2595_),
    .S(_0026_),
    .X(_2869_));
 sky130_fd_sc_hd__buf_1 _5859_ (.A(_2869_),
    .X(_0544_));
 sky130_fd_sc_hd__mux2_2 _5860_ (.A0(\tree_instances[1].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1834_),
    .S(_0026_),
    .X(_2870_));
 sky130_fd_sc_hd__buf_1 _5861_ (.A(_2870_),
    .X(_0545_));
 sky130_fd_sc_hd__mux2_2 _5862_ (.A0(\tree_instances[1].u_tree.pipeline_frame_id[0][4] ),
    .A1(\tree_instances[0].u_tree.frame_id_in[4] ),
    .S(_0026_),
    .X(_2871_));
 sky130_fd_sc_hd__buf_1 _5863_ (.A(_2871_),
    .X(_0546_));
 sky130_fd_sc_hd__inv_2 _5864_ (.A(\tree_instances[1].u_tree.read_enable ),
    .Y(_2872_));
 sky130_fd_sc_hd__buf_1 _5865_ (.A(_2872_),
    .X(_2873_));
 sky130_fd_sc_hd__and2b_2 _5866_ (.A_N(\tree_instances[1].u_tree.tree_state[1] ),
    .B(_2856_),
    .X(_2874_));
 sky130_fd_sc_hd__o21ai_2 _5867_ (.A1(_2873_),
    .A2(_2874_),
    .B1(_2534_),
    .Y(_0547_));
 sky130_fd_sc_hd__mux2_2 _5868_ (.A0(\tree_instances[1].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[1].u_tree.pipeline_frame_id[0][0] ),
    .S(_1227_),
    .X(_2875_));
 sky130_fd_sc_hd__buf_1 _5869_ (.A(_2875_),
    .X(_0548_));
 sky130_fd_sc_hd__mux2_2 _5870_ (.A0(\tree_instances[1].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[1].u_tree.pipeline_frame_id[0][1] ),
    .S(_1227_),
    .X(_2876_));
 sky130_fd_sc_hd__buf_1 _5871_ (.A(_2876_),
    .X(_0549_));
 sky130_fd_sc_hd__mux2_2 _5872_ (.A0(\tree_instances[1].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[1].u_tree.pipeline_frame_id[0][2] ),
    .S(_1227_),
    .X(_2877_));
 sky130_fd_sc_hd__buf_1 _5873_ (.A(_2877_),
    .X(_0550_));
 sky130_fd_sc_hd__mux2_2 _5874_ (.A0(\tree_instances[1].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[1].u_tree.pipeline_frame_id[0][3] ),
    .S(_1227_),
    .X(_2878_));
 sky130_fd_sc_hd__buf_1 _5875_ (.A(_2878_),
    .X(_0551_));
 sky130_fd_sc_hd__mux2_2 _5876_ (.A0(\tree_instances[1].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[1].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[1].u_tree.tree_state[3] ),
    .X(_2879_));
 sky130_fd_sc_hd__buf_1 _5877_ (.A(_2879_),
    .X(_0552_));
 sky130_fd_sc_hd__mux2_2 _5878_ (.A0(\tree_instances[1].u_tree.prediction_out ),
    .A1(\tree_instances[1].u_tree.pipeline_prediction[0][0] ),
    .S(\tree_instances[1].u_tree.tree_state[3] ),
    .X(_2880_));
 sky130_fd_sc_hd__buf_1 _5879_ (.A(_2880_),
    .X(_0553_));
 sky130_fd_sc_hd__a22o_2 _5880_ (.A1(_1227_),
    .A2(_2855_),
    .B1(_1820_),
    .B2(\tree_instances[1].u_tree.ready_for_next ),
    .X(_0554_));
 sky130_fd_sc_hd__inv_2 _5881_ (.A(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .Y(_2881_));
 sky130_fd_sc_hd__inv_2 _5882_ (.A(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .Y(_2882_));
 sky130_fd_sc_hd__a22o_2 _5883_ (.A1(_1404_),
    .A2(_2881_),
    .B1(_2882_),
    .B2(\tree_instances[20].u_tree.pipeline_current_node[0][7] ),
    .X(_2883_));
 sky130_fd_sc_hd__a21o_2 _5884_ (.A1(_1394_),
    .A2(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B1(_2883_),
    .X(_2884_));
 sky130_fd_sc_hd__inv_2 _5885_ (.A(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .Y(_2885_));
 sky130_fd_sc_hd__o221a_2 _5886_ (.A1(_1178_),
    .A2(_2885_),
    .B1(_2882_),
    .B2(\tree_instances[20].u_tree.pipeline_current_node[0][7] ),
    .C1(\tree_instances[20].u_tree.u_tree_weight_rom.cache_valid ),
    .X(_2886_));
 sky130_fd_sc_hd__a22o_2 _5887_ (.A1(_1410_),
    .A2(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .B1(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .B2(_1403_),
    .X(_2887_));
 sky130_fd_sc_hd__a2bb2o_2 _5888_ (.A1_N(_1409_),
    .A2_N(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .B1(_2885_),
    .B2(\tree_instances[20].u_tree.pipeline_current_node[0][5] ),
    .X(_2888_));
 sky130_fd_sc_hd__a221o_2 _5889_ (.A1(_1400_),
    .A2(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .B1(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .B2(_1395_),
    .C1(_2888_),
    .X(_2889_));
 sky130_fd_sc_hd__o22a_2 _5890_ (.A1(_1396_),
    .A2(_2881_),
    .B1(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B2(_1393_),
    .X(_2890_));
 sky130_fd_sc_hd__o221a_2 _5891_ (.A1(_1399_),
    .A2(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .B1(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .B2(_1395_),
    .C1(_2890_),
    .X(_2891_));
 sky130_fd_sc_hd__or2_2 _5892_ (.A(_1403_),
    .B(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .X(_2892_));
 sky130_fd_sc_hd__and4bb_2 _5893_ (.A_N(_2887_),
    .B_N(_2889_),
    .C(_2891_),
    .D(_2892_),
    .X(_2893_));
 sky130_fd_sc_hd__and3b_2 _5894_ (.A_N(_2884_),
    .B(_2886_),
    .C(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__and2b_2 _5895_ (.A_N(_2894_),
    .B(\tree_instances[20].u_tree.read_enable ),
    .X(_2895_));
 sky130_fd_sc_hd__buf_1 _5896_ (.A(_2895_),
    .X(_2896_));
 sky130_fd_sc_hd__buf_1 _5897_ (.A(_2896_),
    .X(_2897_));
 sky130_fd_sc_hd__mux2_2 _5898_ (.A0(\tree_instances[20].u_tree.u_tree_weight_rom.cached_data[12] ),
    .A1(\tree_instances[20].u_tree.u_tree_weight_rom.gen_tree_20.u_tree_rom.node_data[12] ),
    .S(_2897_),
    .X(_2898_));
 sky130_fd_sc_hd__buf_1 _5899_ (.A(_2898_),
    .X(_0555_));
 sky130_fd_sc_hd__buf_1 _5900_ (.A(_2896_),
    .X(_2899_));
 sky130_fd_sc_hd__or3_2 _5901_ (.A(\tree_instances[2].u_tree.tree_state[2] ),
    .B(\tree_instances[2].u_tree.tree_state[1] ),
    .C(_1804_),
    .X(_2900_));
 sky130_fd_sc_hd__buf_1 _5902_ (.A(_2900_),
    .X(_2901_));
 sky130_fd_sc_hd__and2_2 _5903_ (.A(_2147_),
    .B(_2901_),
    .X(_2902_));
 sky130_fd_sc_hd__buf_1 _5904_ (.A(_2902_),
    .X(_0556_));
 sky130_fd_sc_hd__and2_2 _5905_ (.A(_2149_),
    .B(_2901_),
    .X(_2903_));
 sky130_fd_sc_hd__buf_1 _5906_ (.A(_2903_),
    .X(_0557_));
 sky130_fd_sc_hd__and2_2 _5907_ (.A(_2161_),
    .B(_2901_),
    .X(_2904_));
 sky130_fd_sc_hd__buf_1 _5908_ (.A(_2904_),
    .X(_0558_));
 sky130_fd_sc_hd__and2_2 _5909_ (.A(_2163_),
    .B(_2901_),
    .X(_2905_));
 sky130_fd_sc_hd__buf_1 _5910_ (.A(_2905_),
    .X(_0559_));
 sky130_fd_sc_hd__and2_2 _5911_ (.A(_2162_),
    .B(_2901_),
    .X(_2906_));
 sky130_fd_sc_hd__buf_1 _5912_ (.A(_2906_),
    .X(_0560_));
 sky130_fd_sc_hd__and2_2 _5913_ (.A(_2160_),
    .B(_2901_),
    .X(_2907_));
 sky130_fd_sc_hd__buf_1 _5914_ (.A(_2907_),
    .X(_0561_));
 sky130_fd_sc_hd__and2_2 _5915_ (.A(_2157_),
    .B(_2901_),
    .X(_2908_));
 sky130_fd_sc_hd__buf_1 _5916_ (.A(_2908_),
    .X(_0562_));
 sky130_fd_sc_hd__and2_2 _5917_ (.A(_2159_),
    .B(_2900_),
    .X(_2909_));
 sky130_fd_sc_hd__buf_1 _5918_ (.A(_2909_),
    .X(_0563_));
 sky130_fd_sc_hd__and2_2 _5919_ (.A(_2152_),
    .B(_2900_),
    .X(_2910_));
 sky130_fd_sc_hd__buf_1 _5920_ (.A(_2910_),
    .X(_0564_));
 sky130_fd_sc_hd__and2_2 _5921_ (.A(\tree_instances[2].u_tree.pipeline_current_node[0][9] ),
    .B(_2900_),
    .X(_2911_));
 sky130_fd_sc_hd__buf_1 _5922_ (.A(_2911_),
    .X(_0565_));
 sky130_fd_sc_hd__mux2_2 _5923_ (.A0(\tree_instances[2].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1826_),
    .S(_0030_),
    .X(_2912_));
 sky130_fd_sc_hd__buf_1 _5924_ (.A(_2912_),
    .X(_0566_));
 sky130_fd_sc_hd__mux2_2 _5925_ (.A0(\tree_instances[2].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1829_),
    .S(_0030_),
    .X(_2913_));
 sky130_fd_sc_hd__buf_1 _5926_ (.A(_2913_),
    .X(_0567_));
 sky130_fd_sc_hd__mux2_2 _5927_ (.A0(\tree_instances[2].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2595_),
    .S(_0030_),
    .X(_2914_));
 sky130_fd_sc_hd__buf_1 _5928_ (.A(_2914_),
    .X(_0568_));
 sky130_fd_sc_hd__mux2_2 _5929_ (.A0(\tree_instances[2].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1834_),
    .S(_0030_),
    .X(_2915_));
 sky130_fd_sc_hd__buf_1 _5930_ (.A(_2915_),
    .X(_0569_));
 sky130_fd_sc_hd__mux2_2 _5931_ (.A0(\tree_instances[2].u_tree.pipeline_frame_id[0][4] ),
    .A1(\tree_instances[0].u_tree.frame_id_in[4] ),
    .S(_0030_),
    .X(_2916_));
 sky130_fd_sc_hd__buf_1 _5932_ (.A(_2916_),
    .X(_0570_));
 sky130_fd_sc_hd__mux2_2 _5933_ (.A0(\tree_instances[20].u_tree.current_node_data[12] ),
    .A1(\tree_instances[20].u_tree.node_data[12] ),
    .S(_0757_),
    .X(_2917_));
 sky130_fd_sc_hd__buf_1 _5934_ (.A(_2917_),
    .X(_0571_));
 sky130_fd_sc_hd__mux2_2 _5935_ (.A0(\tree_instances[2].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[2].u_tree.pipeline_frame_id[0][0] ),
    .S(_0755_),
    .X(_2918_));
 sky130_fd_sc_hd__buf_1 _5936_ (.A(_2918_),
    .X(_0572_));
 sky130_fd_sc_hd__mux2_2 _5937_ (.A0(\tree_instances[2].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[2].u_tree.pipeline_frame_id[0][1] ),
    .S(_0755_),
    .X(_2919_));
 sky130_fd_sc_hd__buf_1 _5938_ (.A(_2919_),
    .X(_0573_));
 sky130_fd_sc_hd__mux2_2 _5939_ (.A0(\tree_instances[2].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[2].u_tree.pipeline_frame_id[0][2] ),
    .S(_0755_),
    .X(_2920_));
 sky130_fd_sc_hd__buf_1 _5940_ (.A(_2920_),
    .X(_0574_));
 sky130_fd_sc_hd__mux2_2 _5941_ (.A0(\tree_instances[2].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[2].u_tree.pipeline_frame_id[0][3] ),
    .S(_0755_),
    .X(_2921_));
 sky130_fd_sc_hd__buf_1 _5942_ (.A(_2921_),
    .X(_0575_));
 sky130_fd_sc_hd__mux2_2 _5943_ (.A0(\tree_instances[2].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[2].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[2].u_tree.tree_state[3] ),
    .X(_2922_));
 sky130_fd_sc_hd__buf_1 _5944_ (.A(_2922_),
    .X(_0576_));
 sky130_fd_sc_hd__and2_2 _5945_ (.A(_1407_),
    .B(_2553_),
    .X(_2923_));
 sky130_fd_sc_hd__buf_1 _5946_ (.A(_2923_),
    .X(_0577_));
 sky130_fd_sc_hd__and2_2 _5947_ (.A(_1422_),
    .B(_2553_),
    .X(_2924_));
 sky130_fd_sc_hd__buf_1 _5948_ (.A(_2924_),
    .X(_0578_));
 sky130_fd_sc_hd__and2_2 _5949_ (.A(_1431_),
    .B(_2553_),
    .X(_2925_));
 sky130_fd_sc_hd__buf_1 _5950_ (.A(_2925_),
    .X(_0579_));
 sky130_fd_sc_hd__and2_2 _5951_ (.A(_1432_),
    .B(_2553_),
    .X(_2926_));
 sky130_fd_sc_hd__buf_1 _5952_ (.A(_2926_),
    .X(_0580_));
 sky130_fd_sc_hd__and2_2 _5953_ (.A(_1421_),
    .B(_2553_),
    .X(_2927_));
 sky130_fd_sc_hd__buf_1 _5954_ (.A(_2927_),
    .X(_0581_));
 sky130_fd_sc_hd__and2_2 _5955_ (.A(_1424_),
    .B(_2553_),
    .X(_2928_));
 sky130_fd_sc_hd__buf_1 _5956_ (.A(_2928_),
    .X(_0582_));
 sky130_fd_sc_hd__and2_2 _5957_ (.A(_1433_),
    .B(_2553_),
    .X(_2929_));
 sky130_fd_sc_hd__buf_1 _5958_ (.A(_2929_),
    .X(_0583_));
 sky130_fd_sc_hd__and2_2 _5959_ (.A(_1418_),
    .B(_2552_),
    .X(_2930_));
 sky130_fd_sc_hd__buf_1 _5960_ (.A(_2930_),
    .X(_0584_));
 sky130_fd_sc_hd__a22o_2 _5961_ (.A1(_0755_),
    .A2(_2570_),
    .B1(_1804_),
    .B2(\tree_instances[2].u_tree.ready_for_next ),
    .X(_0585_));
 sky130_fd_sc_hd__nand2_2 _5962_ (.A(\tree_instances[7].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[7].u_tree.tree_state[0] ),
    .Y(_2931_));
 sky130_fd_sc_hd__o2bb2a_2 _5963_ (.A1_N(_0970_),
    .A2_N(_2931_),
    .B1(_0040_),
    .B2(\tree_instances[7].u_tree.pipeline_valid[0] ),
    .X(_0586_));
 sky130_fd_sc_hd__buf_1 _5964_ (.A(_0850_),
    .X(_2932_));
 sky130_fd_sc_hd__a22o_2 _5965_ (.A1(\tree_instances[3].u_tree.tree_state[1] ),
    .A2(\tree_instances[3].u_tree.current_node_data[107] ),
    .B1(\tree_instances[3].u_tree.node_data[107] ),
    .B2(_2932_),
    .X(_2933_));
 sky130_fd_sc_hd__o31ai_2 _5966_ (.A1(\tree_instances[3].u_tree.tree_state[0] ),
    .A2(_0850_),
    .A3(\tree_instances[3].u_tree.tree_state[1] ),
    .B1(_0800_),
    .Y(_2934_));
 sky130_fd_sc_hd__nor2_2 _5967_ (.A(_0031_),
    .B(_2934_),
    .Y(_2935_));
 sky130_fd_sc_hd__mux2_2 _5968_ (.A0(\tree_instances[3].u_tree.pipeline_prediction[0][0] ),
    .A1(_2933_),
    .S(_2935_),
    .X(_2936_));
 sky130_fd_sc_hd__buf_1 _5969_ (.A(_2936_),
    .X(_0587_));
 sky130_fd_sc_hd__xor2_2 _5970_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][7] ),
    .B(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .X(_2937_));
 sky130_fd_sc_hd__xor2_2 _5971_ (.A(_1323_),
    .B(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .X(_2938_));
 sky130_fd_sc_hd__inv_2 _5972_ (.A(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .Y(_2939_));
 sky130_fd_sc_hd__a22o_2 _5973_ (.A1(_1328_),
    .A2(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .B1(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B2(_1335_),
    .X(_2940_));
 sky130_fd_sc_hd__xor2_2 _5974_ (.A(\tree_instances[3].u_tree.pipeline_current_node[0][5] ),
    .B(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .X(_2941_));
 sky130_fd_sc_hd__a221o_2 _5975_ (.A1(_1322_),
    .A2(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .B1(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .B2(_1319_),
    .C1(_2941_),
    .X(_2942_));
 sky130_fd_sc_hd__a211o_2 _5976_ (.A1(_1189_),
    .A2(_2939_),
    .B1(_2940_),
    .C1(_2942_),
    .X(_2943_));
 sky130_fd_sc_hd__o22a_2 _5977_ (.A1(_1329_),
    .A2(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .B1(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .B2(_1319_),
    .X(_2944_));
 sky130_fd_sc_hd__o221a_2 _5978_ (.A1(\tree_instances[3].u_tree.pipeline_current_node[0][0] ),
    .A2(_2939_),
    .B1(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .B2(_1322_),
    .C1(\tree_instances[3].u_tree.u_tree_weight_rom.cache_valid ),
    .X(_2945_));
 sky130_fd_sc_hd__o211a_2 _5979_ (.A1(_1335_),
    .A2(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B1(_2944_),
    .C1(_2945_),
    .X(_2946_));
 sky130_fd_sc_hd__or4b_2 _5980_ (.A(_2937_),
    .B(_2938_),
    .C(_2943_),
    .D_N(_2946_),
    .X(_2947_));
 sky130_fd_sc_hd__and2_2 _5981_ (.A(\tree_instances[3].u_tree.read_enable ),
    .B(_2947_),
    .X(_2948_));
 sky130_fd_sc_hd__buf_1 _5982_ (.A(_2948_),
    .X(_2949_));
 sky130_fd_sc_hd__buf_1 _5983_ (.A(_2949_),
    .X(_2950_));
 sky130_fd_sc_hd__buf_1 _5984_ (.A(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__or2_2 _5985_ (.A(\tree_instances[3].u_tree.u_tree_weight_rom.cache_valid ),
    .B(_2951_),
    .X(_2952_));
 sky130_fd_sc_hd__buf_1 _5986_ (.A(_2952_),
    .X(_0588_));
 sky130_fd_sc_hd__mux2_2 _5987_ (.A0(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .A1(_1407_),
    .S(_2899_),
    .X(_2953_));
 sky130_fd_sc_hd__buf_1 _5988_ (.A(_2953_),
    .X(_0589_));
 sky130_fd_sc_hd__mux2_2 _5989_ (.A0(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .A1(_1422_),
    .S(_2899_),
    .X(_2954_));
 sky130_fd_sc_hd__buf_1 _5990_ (.A(_2954_),
    .X(_0590_));
 sky130_fd_sc_hd__mux2_2 _5991_ (.A0(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .A1(_1431_),
    .S(_2899_),
    .X(_2955_));
 sky130_fd_sc_hd__buf_1 _5992_ (.A(_2955_),
    .X(_0591_));
 sky130_fd_sc_hd__mux2_2 _5993_ (.A0(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .A1(_1432_),
    .S(_2899_),
    .X(_2956_));
 sky130_fd_sc_hd__buf_1 _5994_ (.A(_2956_),
    .X(_0592_));
 sky130_fd_sc_hd__mux2_2 _5995_ (.A0(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .A1(_1421_),
    .S(_2899_),
    .X(_2957_));
 sky130_fd_sc_hd__buf_1 _5996_ (.A(_2957_),
    .X(_0593_));
 sky130_fd_sc_hd__mux2_2 _5997_ (.A0(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .A1(_1424_),
    .S(_2899_),
    .X(_2958_));
 sky130_fd_sc_hd__buf_1 _5998_ (.A(_2958_),
    .X(_0594_));
 sky130_fd_sc_hd__buf_1 _5999_ (.A(_2895_),
    .X(_2959_));
 sky130_fd_sc_hd__mux2_2 _6000_ (.A0(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .A1(_1428_),
    .S(_2959_),
    .X(_2960_));
 sky130_fd_sc_hd__buf_1 _6001_ (.A(_2960_),
    .X(_0595_));
 sky130_fd_sc_hd__mux2_2 _6002_ (.A0(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .A1(_1425_),
    .S(_2959_),
    .X(_2961_));
 sky130_fd_sc_hd__buf_1 _6003_ (.A(_2961_),
    .X(_0596_));
 sky130_fd_sc_hd__mux2_2 _6004_ (.A0(\tree_instances[3].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1826_),
    .S(_0032_),
    .X(_2962_));
 sky130_fd_sc_hd__buf_1 _6005_ (.A(_2962_),
    .X(_0597_));
 sky130_fd_sc_hd__mux2_2 _6006_ (.A0(\tree_instances[3].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1829_),
    .S(_0032_),
    .X(_2963_));
 sky130_fd_sc_hd__buf_1 _6007_ (.A(_2963_),
    .X(_0598_));
 sky130_fd_sc_hd__mux2_2 _6008_ (.A0(\tree_instances[3].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2595_),
    .S(_0032_),
    .X(_2964_));
 sky130_fd_sc_hd__buf_1 _6009_ (.A(_2964_),
    .X(_0599_));
 sky130_fd_sc_hd__mux2_2 _6010_ (.A0(\tree_instances[3].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1834_),
    .S(_0032_),
    .X(_2965_));
 sky130_fd_sc_hd__buf_1 _6011_ (.A(_2965_),
    .X(_0600_));
 sky130_fd_sc_hd__mux2_2 _6012_ (.A0(\tree_instances[3].u_tree.pipeline_frame_id[0][4] ),
    .A1(\tree_instances[0].u_tree.frame_id_in[4] ),
    .S(_0032_),
    .X(_2966_));
 sky130_fd_sc_hd__buf_1 _6013_ (.A(_2966_),
    .X(_0601_));
 sky130_fd_sc_hd__inv_2 _6014_ (.A(_0032_),
    .Y(_2967_));
 sky130_fd_sc_hd__inv_2 _6015_ (.A(\tree_instances[3].u_tree.read_enable ),
    .Y(_2968_));
 sky130_fd_sc_hd__buf_1 _6016_ (.A(_2968_),
    .X(_2969_));
 sky130_fd_sc_hd__o21ba_2 _6017_ (.A1(\tree_instances[3].u_tree.tree_state[0] ),
    .A2(_0851_),
    .B1_N(\tree_instances[3].u_tree.tree_state[1] ),
    .X(_2970_));
 sky130_fd_sc_hd__or3_2 _6018_ (.A(\tree_instances[3].u_tree.tree_state[2] ),
    .B(\tree_instances[3].u_tree.tree_state[1] ),
    .C(_2967_),
    .X(_2971_));
 sky130_fd_sc_hd__buf_1 _6019_ (.A(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__o21ai_2 _6020_ (.A1(_2969_),
    .A2(_2970_),
    .B1(_2972_),
    .Y(_0602_));
 sky130_fd_sc_hd__mux2_2 _6021_ (.A0(\tree_instances[3].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[3].u_tree.pipeline_frame_id[0][0] ),
    .S(_0799_),
    .X(_2973_));
 sky130_fd_sc_hd__buf_1 _6022_ (.A(_2973_),
    .X(_0603_));
 sky130_fd_sc_hd__mux2_2 _6023_ (.A0(\tree_instances[3].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[3].u_tree.pipeline_frame_id[0][1] ),
    .S(_0799_),
    .X(_2974_));
 sky130_fd_sc_hd__buf_1 _6024_ (.A(_2974_),
    .X(_0604_));
 sky130_fd_sc_hd__mux2_2 _6025_ (.A0(\tree_instances[3].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[3].u_tree.pipeline_frame_id[0][2] ),
    .S(_0799_),
    .X(_2975_));
 sky130_fd_sc_hd__buf_1 _6026_ (.A(_2975_),
    .X(_0605_));
 sky130_fd_sc_hd__mux2_2 _6027_ (.A0(\tree_instances[3].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[3].u_tree.pipeline_frame_id[0][3] ),
    .S(_0799_),
    .X(_2976_));
 sky130_fd_sc_hd__buf_1 _6028_ (.A(_2976_),
    .X(_0606_));
 sky130_fd_sc_hd__mux2_2 _6029_ (.A0(\tree_instances[3].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[3].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[3].u_tree.tree_state[3] ),
    .X(_2977_));
 sky130_fd_sc_hd__buf_1 _6030_ (.A(_2977_),
    .X(_0607_));
 sky130_fd_sc_hd__mux2_2 _6031_ (.A0(\tree_instances[3].u_tree.prediction_out ),
    .A1(\tree_instances[3].u_tree.pipeline_prediction[0][0] ),
    .S(\tree_instances[3].u_tree.tree_state[3] ),
    .X(_2978_));
 sky130_fd_sc_hd__buf_1 _6032_ (.A(_2978_),
    .X(_0608_));
 sky130_fd_sc_hd__a22o_2 _6033_ (.A1(_0799_),
    .A2(_0800_),
    .B1(_2967_),
    .B2(\tree_instances[3].u_tree.ready_for_next ),
    .X(_0609_));
 sky130_fd_sc_hd__nor2_2 _6034_ (.A(_2872_),
    .B(_2517_),
    .Y(_2979_));
 sky130_fd_sc_hd__buf_1 _6035_ (.A(_2979_),
    .X(_2980_));
 sky130_fd_sc_hd__buf_1 _6036_ (.A(_2980_),
    .X(_2981_));
 sky130_fd_sc_hd__a221o_2 _6037_ (.A1(_2873_),
    .A2(\tree_instances[1].u_tree.node_data[12] ),
    .B1(\tree_instances[1].u_tree.u_tree_weight_rom.cached_data[12] ),
    .B2(_2981_),
    .C1(_2532_),
    .X(_0610_));
 sky130_fd_sc_hd__nor2_2 _6038_ (.A(_2968_),
    .B(_2947_),
    .Y(_2982_));
 sky130_fd_sc_hd__buf_1 _6039_ (.A(_2982_),
    .X(_2983_));
 sky130_fd_sc_hd__buf_1 _6040_ (.A(_2949_),
    .X(_2984_));
 sky130_fd_sc_hd__buf_1 _6041_ (.A(_2969_),
    .X(_2985_));
 sky130_fd_sc_hd__buf_1 _6042_ (.A(_2983_),
    .X(_2986_));
 sky130_fd_sc_hd__a22o_2 _6043_ (.A1(\tree_instances[3].u_tree.u_tree_weight_rom.gen_tree_3.u_tree_rom.node_data[107] ),
    .A2(_2984_),
    .B1(_2986_),
    .B2(\tree_instances[3].u_tree.u_tree_weight_rom.cached_data[107] ),
    .X(_2987_));
 sky130_fd_sc_hd__a21o_2 _6044_ (.A1(_2985_),
    .A2(\tree_instances[3].u_tree.node_data[107] ),
    .B1(_2987_),
    .X(_0611_));
 sky130_fd_sc_hd__buf_1 _6045_ (.A(_2949_),
    .X(_2988_));
 sky130_fd_sc_hd__buf_1 _6046_ (.A(_2988_),
    .X(_2989_));
 sky130_fd_sc_hd__and2_2 _6047_ (.A(_2452_),
    .B(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .X(_2990_));
 sky130_fd_sc_hd__nor2_2 _6048_ (.A(_0937_),
    .B(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .Y(_2991_));
 sky130_fd_sc_hd__o221a_2 _6049_ (.A1(_2450_),
    .A2(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .B1(_2990_),
    .B2(_2991_),
    .C1(\tree_instances[5].u_tree.u_tree_weight_rom.cache_valid ),
    .X(_2992_));
 sky130_fd_sc_hd__inv_2 _6050_ (.A(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .Y(_2993_));
 sky130_fd_sc_hd__a22o_2 _6051_ (.A1(_1247_),
    .A2(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B1(_2993_),
    .B2(\tree_instances[5].u_tree.pipeline_current_node[0][7] ),
    .X(_2994_));
 sky130_fd_sc_hd__a221oi_2 _6052_ (.A1(_2450_),
    .A2(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .B1(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .B2(_2465_),
    .C1(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__inv_2 _6053_ (.A(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .Y(_2996_));
 sky130_fd_sc_hd__o22a_2 _6054_ (.A1(_1247_),
    .A2(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .B1(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[8] ),
    .B2(_2472_),
    .X(_2997_));
 sky130_fd_sc_hd__inv_2 _6055_ (.A(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[8] ),
    .Y(_2998_));
 sky130_fd_sc_hd__o2bb2a_2 _6056_ (.A1_N(_2464_),
    .A2_N(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .B1(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .B2(_2460_),
    .X(_2999_));
 sky130_fd_sc_hd__o221a_2 _6057_ (.A1(\tree_instances[5].u_tree.pipeline_current_node[0][7] ),
    .A2(_2993_),
    .B1(_2998_),
    .B2(\tree_instances[5].u_tree.pipeline_current_node[0][8] ),
    .C1(_2999_),
    .X(_3000_));
 sky130_fd_sc_hd__xnor2_2 _6058_ (.A(\tree_instances[5].u_tree.pipeline_current_node[0][4] ),
    .B(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .Y(_3001_));
 sky130_fd_sc_hd__o221a_2 _6059_ (.A1(_2465_),
    .A2(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .B1(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .B2(_2464_),
    .C1(_3001_),
    .X(_3002_));
 sky130_fd_sc_hd__o2111a_2 _6060_ (.A1(_1240_),
    .A2(_2996_),
    .B1(_2997_),
    .C1(_3000_),
    .D1(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__inv_2 _6061_ (.A(\tree_instances[5].u_tree.read_enable ),
    .Y(_3004_));
 sky130_fd_sc_hd__a31o_2 _6062_ (.A1(_2992_),
    .A2(_2995_),
    .A3(_3003_),
    .B1(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__and4_2 _6063_ (.A(_1248_),
    .B(_2483_),
    .C(_2485_),
    .D(_2492_),
    .X(_3006_));
 sky130_fd_sc_hd__a2111oi_2 _6064_ (.A1(\tree_instances[5].u_tree.pipeline_current_node[0][7] ),
    .A2(_2489_),
    .B1(_3005_),
    .C1(_3006_),
    .D1(\tree_instances[5].u_tree.pipeline_current_node[0][8] ),
    .Y(_3007_));
 sky130_fd_sc_hd__buf_1 _6065_ (.A(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__buf_1 _6066_ (.A(_3008_),
    .X(_3009_));
 sky130_fd_sc_hd__buf_1 _6067_ (.A(_3009_),
    .X(_3010_));
 sky130_fd_sc_hd__buf_1 _6068_ (.A(_3005_),
    .X(_3011_));
 sky130_fd_sc_hd__buf_1 _6069_ (.A(_3009_),
    .X(_3012_));
 sky130_fd_sc_hd__buf_1 _6070_ (.A(_3005_),
    .X(_3013_));
 sky130_fd_sc_hd__buf_1 _6071_ (.A(\tree_instances[5].u_tree.read_enable ),
    .X(_3014_));
 sky130_fd_sc_hd__mux2_2 _6072_ (.A0(\tree_instances[5].u_tree.node_data[107] ),
    .A1(\tree_instances[5].u_tree.u_tree_weight_rom.cached_data[107] ),
    .S(_3014_),
    .X(_3015_));
 sky130_fd_sc_hd__a22o_2 _6073_ (.A1(\tree_instances[5].u_tree.u_tree_weight_rom.gen_tree_5.u_tree_rom.node_data[107] ),
    .A2(_3012_),
    .B1(_3015_),
    .B2(_3013_),
    .X(_0612_));
 sky130_fd_sc_hd__mux2_2 _6074_ (.A0(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .A1(_1325_),
    .S(_2989_),
    .X(_3016_));
 sky130_fd_sc_hd__buf_1 _6075_ (.A(_3016_),
    .X(_0613_));
 sky130_fd_sc_hd__mux2_2 _6076_ (.A0(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .A1(_1351_),
    .S(_2989_),
    .X(_3017_));
 sky130_fd_sc_hd__buf_1 _6077_ (.A(_3017_),
    .X(_0614_));
 sky130_fd_sc_hd__mux2_2 _6078_ (.A0(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .A1(_1350_),
    .S(_2989_),
    .X(_3018_));
 sky130_fd_sc_hd__buf_1 _6079_ (.A(_3018_),
    .X(_0615_));
 sky130_fd_sc_hd__mux2_2 _6080_ (.A0(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .A1(_1347_),
    .S(_2989_),
    .X(_3019_));
 sky130_fd_sc_hd__buf_1 _6081_ (.A(_3019_),
    .X(_0616_));
 sky130_fd_sc_hd__buf_1 _6082_ (.A(_2988_),
    .X(_3020_));
 sky130_fd_sc_hd__mux2_2 _6083_ (.A0(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .A1(_1344_),
    .S(_3020_),
    .X(_3021_));
 sky130_fd_sc_hd__buf_1 _6084_ (.A(_3021_),
    .X(_0617_));
 sky130_fd_sc_hd__mux2_2 _6085_ (.A0(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .A1(_1352_),
    .S(_3020_),
    .X(_3022_));
 sky130_fd_sc_hd__buf_1 _6086_ (.A(_3022_),
    .X(_0618_));
 sky130_fd_sc_hd__mux2_2 _6087_ (.A0(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .A1(_1327_),
    .S(_3020_),
    .X(_3023_));
 sky130_fd_sc_hd__buf_1 _6088_ (.A(_3023_),
    .X(_0619_));
 sky130_fd_sc_hd__mux2_2 _6089_ (.A0(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .A1(_1346_),
    .S(_3020_),
    .X(_3024_));
 sky130_fd_sc_hd__buf_1 _6090_ (.A(_3024_),
    .X(_0620_));
 sky130_fd_sc_hd__buf_1 _6091_ (.A(_2988_),
    .X(_3025_));
 sky130_fd_sc_hd__mux2_2 _6092_ (.A0(\tree_instances[3].u_tree.u_tree_weight_rom.cached_data[107] ),
    .A1(\tree_instances[3].u_tree.u_tree_weight_rom.gen_tree_3.u_tree_rom.node_data[107] ),
    .S(_3025_),
    .X(_3026_));
 sky130_fd_sc_hd__buf_1 _6093_ (.A(_3026_),
    .X(_0621_));
 sky130_fd_sc_hd__mux2_2 _6094_ (.A0(\tree_instances[4].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1826_),
    .S(_0034_),
    .X(_3027_));
 sky130_fd_sc_hd__buf_1 _6095_ (.A(_3027_),
    .X(_0622_));
 sky130_fd_sc_hd__mux2_2 _6096_ (.A0(\tree_instances[4].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1829_),
    .S(_0034_),
    .X(_3028_));
 sky130_fd_sc_hd__buf_1 _6097_ (.A(_3028_),
    .X(_0623_));
 sky130_fd_sc_hd__mux2_2 _6098_ (.A0(\tree_instances[4].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2595_),
    .S(_0034_),
    .X(_3029_));
 sky130_fd_sc_hd__buf_1 _6099_ (.A(_3029_),
    .X(_0624_));
 sky130_fd_sc_hd__mux2_2 _6100_ (.A0(\tree_instances[4].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1834_),
    .S(_0034_),
    .X(_3030_));
 sky130_fd_sc_hd__buf_1 _6101_ (.A(_3030_),
    .X(_0625_));
 sky130_fd_sc_hd__mux2_2 _6102_ (.A0(\tree_instances[4].u_tree.pipeline_frame_id[0][4] ),
    .A1(\tree_instances[0].u_tree.frame_id_in[4] ),
    .S(_0034_),
    .X(_3031_));
 sky130_fd_sc_hd__buf_1 _6103_ (.A(_3031_),
    .X(_0626_));
 sky130_fd_sc_hd__buf_1 _6104_ (.A(_2932_),
    .X(_3032_));
 sky130_fd_sc_hd__mux2_2 _6105_ (.A0(\tree_instances[3].u_tree.current_node_data[107] ),
    .A1(\tree_instances[3].u_tree.node_data[107] ),
    .S(_3032_),
    .X(_3033_));
 sky130_fd_sc_hd__buf_1 _6106_ (.A(_3033_),
    .X(_0627_));
 sky130_fd_sc_hd__or3_2 _6107_ (.A(\tree_instances[4].u_tree.tree_state[1] ),
    .B(\tree_instances[4].u_tree.tree_state[2] ),
    .C(_1807_),
    .X(_3034_));
 sky130_fd_sc_hd__buf_1 _6108_ (.A(_3034_),
    .X(_3035_));
 sky130_fd_sc_hd__mux2_2 _6109_ (.A0(\tree_instances[4].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[4].u_tree.pipeline_frame_id[0][0] ),
    .S(_0849_),
    .X(_3036_));
 sky130_fd_sc_hd__buf_1 _6110_ (.A(_3036_),
    .X(_0628_));
 sky130_fd_sc_hd__mux2_2 _6111_ (.A0(\tree_instances[4].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[4].u_tree.pipeline_frame_id[0][1] ),
    .S(_0849_),
    .X(_3037_));
 sky130_fd_sc_hd__buf_1 _6112_ (.A(_3037_),
    .X(_0629_));
 sky130_fd_sc_hd__mux2_2 _6113_ (.A0(\tree_instances[4].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[4].u_tree.pipeline_frame_id[0][2] ),
    .S(_0849_),
    .X(_3038_));
 sky130_fd_sc_hd__buf_1 _6114_ (.A(_3038_),
    .X(_0630_));
 sky130_fd_sc_hd__mux2_2 _6115_ (.A0(\tree_instances[4].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[4].u_tree.pipeline_frame_id[0][3] ),
    .S(_0849_),
    .X(_3039_));
 sky130_fd_sc_hd__buf_1 _6116_ (.A(_3039_),
    .X(_0631_));
 sky130_fd_sc_hd__mux2_2 _6117_ (.A0(\tree_instances[4].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[4].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[4].u_tree.tree_state[3] ),
    .X(_3040_));
 sky130_fd_sc_hd__buf_1 _6118_ (.A(_3040_),
    .X(_0632_));
 sky130_fd_sc_hd__and2_2 _6119_ (.A(_1325_),
    .B(_2972_),
    .X(_3041_));
 sky130_fd_sc_hd__buf_1 _6120_ (.A(_3041_),
    .X(_0633_));
 sky130_fd_sc_hd__and2_2 _6121_ (.A(_1351_),
    .B(_2972_),
    .X(_3042_));
 sky130_fd_sc_hd__buf_1 _6122_ (.A(_3042_),
    .X(_0634_));
 sky130_fd_sc_hd__and2_2 _6123_ (.A(_1350_),
    .B(_2972_),
    .X(_3043_));
 sky130_fd_sc_hd__buf_1 _6124_ (.A(_3043_),
    .X(_0635_));
 sky130_fd_sc_hd__and2_2 _6125_ (.A(_1347_),
    .B(_2972_),
    .X(_3044_));
 sky130_fd_sc_hd__buf_1 _6126_ (.A(_3044_),
    .X(_0636_));
 sky130_fd_sc_hd__and2_2 _6127_ (.A(_1344_),
    .B(_2972_),
    .X(_3045_));
 sky130_fd_sc_hd__buf_1 _6128_ (.A(_3045_),
    .X(_0637_));
 sky130_fd_sc_hd__and2_2 _6129_ (.A(_1352_),
    .B(_2972_),
    .X(_3046_));
 sky130_fd_sc_hd__buf_1 _6130_ (.A(_3046_),
    .X(_0638_));
 sky130_fd_sc_hd__and2_2 _6131_ (.A(_1327_),
    .B(_2972_),
    .X(_3047_));
 sky130_fd_sc_hd__buf_1 _6132_ (.A(_3047_),
    .X(_0639_));
 sky130_fd_sc_hd__and2_2 _6133_ (.A(_1346_),
    .B(_2971_),
    .X(_3048_));
 sky130_fd_sc_hd__buf_1 _6134_ (.A(_3048_),
    .X(_0640_));
 sky130_fd_sc_hd__a22o_2 _6135_ (.A1(_0849_),
    .A2(_1955_),
    .B1(_1807_),
    .B2(\tree_instances[4].u_tree.ready_for_next ),
    .X(_0641_));
 sky130_fd_sc_hd__nand2_2 _6136_ (.A(\tree_instances[17].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[17].u_tree.tree_state[0] ),
    .Y(_3049_));
 sky130_fd_sc_hd__o2bb2a_2 _6137_ (.A1_N(_0909_),
    .A2_N(_3049_),
    .B1(_0020_),
    .B2(\tree_instances[17].u_tree.pipeline_valid[0] ),
    .X(_0642_));
 sky130_fd_sc_hd__buf_1 _6138_ (.A(_2130_),
    .X(_3050_));
 sky130_fd_sc_hd__nand3_2 _6139_ (.A(_2104_),
    .B(_2105_),
    .C(_2106_),
    .Y(_3051_));
 sky130_fd_sc_hd__and4_2 _6140_ (.A(\tree_instances[12].u_tree.u_tree_weight_rom.cache_valid ),
    .B(_2100_),
    .C(_2101_),
    .D(_2102_),
    .X(_3052_));
 sky130_fd_sc_hd__or2b_2 _6141_ (.A(_2099_),
    .B_N(_3052_),
    .X(_3053_));
 sky130_fd_sc_hd__nor4_2 _6142_ (.A(_2129_),
    .B(_2093_),
    .C(_3051_),
    .D(_3053_),
    .Y(_3054_));
 sky130_fd_sc_hd__buf_1 _6143_ (.A(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__a22o_2 _6144_ (.A1(\tree_instances[12].u_tree.u_tree_weight_rom.gen_tree_12.u_tree_rom.node_data[12] ),
    .A2(_2112_),
    .B1(_3055_),
    .B2(\tree_instances[12].u_tree.u_tree_weight_rom.cached_data[12] ),
    .X(_3056_));
 sky130_fd_sc_hd__a21o_2 _6145_ (.A1(_3050_),
    .A2(\tree_instances[12].u_tree.node_data[12] ),
    .B1(_3056_),
    .X(_0643_));
 sky130_fd_sc_hd__nand2_2 _6146_ (.A(_1661_),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .Y(_3057_));
 sky130_fd_sc_hd__or2_2 _6147_ (.A(\tree_instances[13].u_tree.pipeline_current_node[0][6] ),
    .B(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .X(_3058_));
 sky130_fd_sc_hd__a221o_2 _6148_ (.A1(_1686_),
    .A2(_2170_),
    .B1(_3057_),
    .B2(_3058_),
    .C1(_2169_),
    .X(_3059_));
 sky130_fd_sc_hd__or4_2 _6149_ (.A(_2176_),
    .B(_2179_),
    .C(_2183_),
    .D(_2184_),
    .X(_3060_));
 sky130_fd_sc_hd__o21ai_2 _6150_ (.A1(_1658_),
    .A2(_2170_),
    .B1(_2173_),
    .Y(_3061_));
 sky130_fd_sc_hd__or4_2 _6151_ (.A(_3060_),
    .B(_3061_),
    .C(_2178_),
    .D(_2185_),
    .X(_3062_));
 sky130_fd_sc_hd__or4b_2 _6152_ (.A(_2175_),
    .B(_3062_),
    .C(_2182_),
    .D_N(_2172_),
    .X(_3063_));
 sky130_fd_sc_hd__nor4_2 _6153_ (.A(_2218_),
    .B(_2171_),
    .C(_3059_),
    .D(_3063_),
    .Y(_3064_));
 sky130_fd_sc_hd__buf_1 _6154_ (.A(_3064_),
    .X(_3065_));
 sky130_fd_sc_hd__buf_1 _6155_ (.A(_3065_),
    .X(_3066_));
 sky130_fd_sc_hd__a221o_2 _6156_ (.A1(_2219_),
    .A2(\tree_instances[13].u_tree.node_data[12] ),
    .B1(_3066_),
    .B2(\tree_instances[13].u_tree.u_tree_weight_rom.cached_data[12] ),
    .C1(_2244_),
    .X(_0644_));
 sky130_fd_sc_hd__nand2_2 _6157_ (.A(\tree_instances[1].u_tree.tree_state[0] ),
    .B(\tree_instances[1].u_tree.pipeline_valid[0] ),
    .Y(_3067_));
 sky130_fd_sc_hd__o2bb2a_2 _6158_ (.A1_N(_1227_),
    .A2_N(_3067_),
    .B1(_0026_),
    .B2(\tree_instances[1].u_tree.pipeline_valid[0] ),
    .X(_0645_));
 sky130_fd_sc_hd__buf_1 _6159_ (.A(_2959_),
    .X(_3068_));
 sky130_fd_sc_hd__and2_2 _6160_ (.A(\tree_instances[20].u_tree.read_enable ),
    .B(_2894_),
    .X(_3069_));
 sky130_fd_sc_hd__buf_1 _6161_ (.A(_3069_),
    .X(_3070_));
 sky130_fd_sc_hd__buf_1 _6162_ (.A(_3070_),
    .X(_3071_));
 sky130_fd_sc_hd__and2b_2 _6163_ (.A_N(_2502_),
    .B(\tree_instances[20].u_tree.node_data[12] ),
    .X(_3072_));
 sky130_fd_sc_hd__a221o_2 _6164_ (.A1(\tree_instances[20].u_tree.u_tree_weight_rom.gen_tree_20.u_tree_rom.node_data[12] ),
    .A2(_3068_),
    .B1(_3071_),
    .B2(\tree_instances[20].u_tree.u_tree_weight_rom.cached_data[12] ),
    .C1(_3072_),
    .X(_0646_));
 sky130_fd_sc_hd__buf_1 _6165_ (.A(_0717_),
    .X(_3073_));
 sky130_fd_sc_hd__buf_1 _6166_ (.A(_3073_),
    .X(_3074_));
 sky130_fd_sc_hd__buf_1 _6167_ (.A(_3074_),
    .X(_3075_));
 sky130_fd_sc_hd__buf_1 _6168_ (.A(_3075_),
    .X(_3076_));
 sky130_fd_sc_hd__buf_1 _6169_ (.A(_2567_),
    .X(_3077_));
 sky130_fd_sc_hd__buf_1 _6170_ (.A(_3077_),
    .X(_3078_));
 sky130_fd_sc_hd__buf_1 _6171_ (.A(_2561_),
    .X(_3079_));
 sky130_fd_sc_hd__buf_1 _6172_ (.A(_3078_),
    .X(_3080_));
 sky130_fd_sc_hd__nand2_2 _6173_ (.A(\tree_instances[6].u_tree.tree_state[0] ),
    .B(_0931_),
    .Y(_3081_));
 sky130_fd_sc_hd__o2bb2a_2 _6174_ (.A1_N(_0932_),
    .A2_N(_3081_),
    .B1(_0038_),
    .B2(\tree_instances[6].u_tree.pipeline_valid[0] ),
    .X(_0647_));
 sky130_fd_sc_hd__a22o_2 _6175_ (.A1(\tree_instances[5].u_tree.tree_state[1] ),
    .A2(\tree_instances[5].u_tree.current_node_data[107] ),
    .B1(\tree_instances[5].u_tree.node_data[107] ),
    .B2(_0933_),
    .X(_3082_));
 sky130_fd_sc_hd__nor3_2 _6176_ (.A(\tree_instances[5].u_tree.tree_state[0] ),
    .B(\tree_instances[5].u_tree.tree_state[1] ),
    .C(\tree_instances[5].u_tree.tree_state[2] ),
    .Y(_3083_));
 sky130_fd_sc_hd__a211oi_2 _6177_ (.A1(\tree_instances[5].u_tree.tree_state[0] ),
    .A2(_0902_),
    .B1(_0035_),
    .C1(_3083_),
    .Y(_3084_));
 sky130_fd_sc_hd__mux2_2 _6178_ (.A0(\tree_instances[5].u_tree.pipeline_prediction[0][0] ),
    .A1(_3082_),
    .S(_3084_),
    .X(_3085_));
 sky130_fd_sc_hd__buf_1 _6179_ (.A(_3085_),
    .X(_0648_));
 sky130_fd_sc_hd__a21o_2 _6180_ (.A1(\tree_instances[5].u_tree.u_tree_weight_rom.cache_valid ),
    .A2(_3011_),
    .B1(_3010_),
    .X(_0649_));
 sky130_fd_sc_hd__and2_2 _6181_ (.A(_3076_),
    .B(_3035_),
    .X(_3086_));
 sky130_fd_sc_hd__buf_1 _6182_ (.A(_3086_),
    .X(_0650_));
 sky130_fd_sc_hd__and2_2 _6183_ (.A(_1888_),
    .B(_3035_),
    .X(_3087_));
 sky130_fd_sc_hd__buf_1 _6184_ (.A(_3087_),
    .X(_0651_));
 sky130_fd_sc_hd__and2_2 _6185_ (.A(_1885_),
    .B(_3035_),
    .X(_3088_));
 sky130_fd_sc_hd__buf_1 _6186_ (.A(_3088_),
    .X(_0652_));
 sky130_fd_sc_hd__and2_2 _6187_ (.A(_2565_),
    .B(_3035_),
    .X(_3089_));
 sky130_fd_sc_hd__buf_1 _6188_ (.A(_3089_),
    .X(_0653_));
 sky130_fd_sc_hd__and2_2 _6189_ (.A(_3080_),
    .B(_3035_),
    .X(_3090_));
 sky130_fd_sc_hd__buf_1 _6190_ (.A(_3090_),
    .X(_0654_));
 sky130_fd_sc_hd__and2_2 _6191_ (.A(_0709_),
    .B(_3035_),
    .X(_3091_));
 sky130_fd_sc_hd__buf_1 _6192_ (.A(_3091_),
    .X(_0655_));
 sky130_fd_sc_hd__and2_2 _6193_ (.A(_1891_),
    .B(_3035_),
    .X(_3092_));
 sky130_fd_sc_hd__buf_1 _6194_ (.A(_3092_),
    .X(_0656_));
 sky130_fd_sc_hd__and2_2 _6195_ (.A(_2563_),
    .B(_3034_),
    .X(_3093_));
 sky130_fd_sc_hd__buf_1 _6196_ (.A(_3093_),
    .X(_0657_));
 sky130_fd_sc_hd__and2_2 _6197_ (.A(_3079_),
    .B(_3034_),
    .X(_3094_));
 sky130_fd_sc_hd__buf_1 _6198_ (.A(_3094_),
    .X(_0658_));
 sky130_fd_sc_hd__mux2_2 _6199_ (.A0(\tree_instances[5].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1826_),
    .S(_0036_),
    .X(_3095_));
 sky130_fd_sc_hd__buf_1 _6200_ (.A(_3095_),
    .X(_0659_));
 sky130_fd_sc_hd__mux2_2 _6201_ (.A0(\tree_instances[5].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1829_),
    .S(_0036_),
    .X(_3096_));
 sky130_fd_sc_hd__buf_1 _6202_ (.A(_3096_),
    .X(_0660_));
 sky130_fd_sc_hd__mux2_2 _6203_ (.A0(\tree_instances[5].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2595_),
    .S(_0036_),
    .X(_3097_));
 sky130_fd_sc_hd__buf_1 _6204_ (.A(_3097_),
    .X(_0661_));
 sky130_fd_sc_hd__mux2_2 _6205_ (.A0(\tree_instances[5].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1834_),
    .S(_0036_),
    .X(_3098_));
 sky130_fd_sc_hd__buf_1 _6206_ (.A(_3098_),
    .X(_0662_));
 sky130_fd_sc_hd__mux2_2 _6207_ (.A0(\tree_instances[5].u_tree.pipeline_frame_id[0][4] ),
    .A1(\tree_instances[0].u_tree.frame_id_in[4] ),
    .S(_0036_),
    .X(_3099_));
 sky130_fd_sc_hd__buf_1 _6208_ (.A(_3099_),
    .X(_0663_));
 sky130_fd_sc_hd__nor2_2 _6209_ (.A(\tree_instances[5].u_tree.tree_state[1] ),
    .B(_3083_),
    .Y(_3100_));
 sky130_fd_sc_hd__or3_2 _6210_ (.A(\tree_instances[5].u_tree.tree_state[1] ),
    .B(\tree_instances[5].u_tree.tree_state[2] ),
    .C(_1808_),
    .X(_3101_));
 sky130_fd_sc_hd__buf_1 _6211_ (.A(_3101_),
    .X(_3102_));
 sky130_fd_sc_hd__o21ai_2 _6212_ (.A1(_3004_),
    .A2(_3100_),
    .B1(_3102_),
    .Y(_0664_));
 sky130_fd_sc_hd__mux2_2 _6213_ (.A0(\tree_instances[5].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[5].u_tree.pipeline_frame_id[0][0] ),
    .S(_0903_),
    .X(_3103_));
 sky130_fd_sc_hd__buf_1 _6214_ (.A(_3103_),
    .X(_0665_));
 sky130_fd_sc_hd__mux2_2 _6215_ (.A0(\tree_instances[5].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[5].u_tree.pipeline_frame_id[0][1] ),
    .S(_0903_),
    .X(_3104_));
 sky130_fd_sc_hd__buf_1 _6216_ (.A(_3104_),
    .X(_0666_));
 sky130_fd_sc_hd__mux2_2 _6217_ (.A0(\tree_instances[5].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[5].u_tree.pipeline_frame_id[0][2] ),
    .S(_0903_),
    .X(_3105_));
 sky130_fd_sc_hd__buf_1 _6218_ (.A(_3105_),
    .X(_0667_));
 sky130_fd_sc_hd__mux2_2 _6219_ (.A0(\tree_instances[5].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[5].u_tree.pipeline_frame_id[0][3] ),
    .S(_0903_),
    .X(_3106_));
 sky130_fd_sc_hd__buf_1 _6220_ (.A(_3106_),
    .X(_0668_));
 sky130_fd_sc_hd__mux2_2 _6221_ (.A0(\tree_instances[5].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[5].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[5].u_tree.tree_state[3] ),
    .X(_3107_));
 sky130_fd_sc_hd__buf_1 _6222_ (.A(_3107_),
    .X(_0669_));
 sky130_fd_sc_hd__mux2_2 _6223_ (.A0(\tree_instances[5].u_tree.prediction_out ),
    .A1(\tree_instances[5].u_tree.pipeline_prediction[0][0] ),
    .S(\tree_instances[5].u_tree.tree_state[3] ),
    .X(_3108_));
 sky130_fd_sc_hd__buf_1 _6224_ (.A(_3108_),
    .X(_0670_));
 sky130_fd_sc_hd__nand2_2 _6225_ (.A(\tree_instances[5].u_tree.tree_state[0] ),
    .B(_0902_),
    .Y(_3109_));
 sky130_fd_sc_hd__a22o_2 _6226_ (.A1(_0903_),
    .A2(_3109_),
    .B1(_1808_),
    .B2(\tree_instances[5].u_tree.ready_for_next ),
    .X(_0671_));
 sky130_fd_sc_hd__buf_1 _6227_ (.A(_2311_),
    .X(_3110_));
 sky130_fd_sc_hd__buf_1 _6228_ (.A(_2361_),
    .X(_3111_));
 sky130_fd_sc_hd__nor2_2 _6229_ (.A(_2310_),
    .B(_2360_),
    .Y(_3112_));
 sky130_fd_sc_hd__buf_1 _6230_ (.A(_3112_),
    .X(_3113_));
 sky130_fd_sc_hd__buf_1 _6231_ (.A(_3113_),
    .X(_3114_));
 sky130_fd_sc_hd__a22o_2 _6232_ (.A1(\tree_instances[16].u_tree.u_tree_weight_rom.gen_tree_16.u_tree_rom.node_data[12] ),
    .A2(_3111_),
    .B1(_3114_),
    .B2(\tree_instances[16].u_tree.u_tree_weight_rom.cached_data[12] ),
    .X(_3115_));
 sky130_fd_sc_hd__a21o_2 _6233_ (.A1(_3110_),
    .A2(\tree_instances[16].u_tree.node_data[12] ),
    .B1(_3115_),
    .X(_0672_));
 sky130_fd_sc_hd__buf_1 _6234_ (.A(_3007_),
    .X(_3116_));
 sky130_fd_sc_hd__mux2_2 _6235_ (.A0(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[0] ),
    .A1(_2456_),
    .S(_3116_),
    .X(_3117_));
 sky130_fd_sc_hd__buf_1 _6236_ (.A(_3117_),
    .X(_0673_));
 sky130_fd_sc_hd__mux2_2 _6237_ (.A0(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[1] ),
    .A1(_2486_),
    .S(_3116_),
    .X(_3118_));
 sky130_fd_sc_hd__buf_1 _6238_ (.A(_3118_),
    .X(_0674_));
 sky130_fd_sc_hd__mux2_2 _6239_ (.A0(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[2] ),
    .A1(_2481_),
    .S(_3116_),
    .X(_3119_));
 sky130_fd_sc_hd__buf_1 _6240_ (.A(_3119_),
    .X(_0675_));
 sky130_fd_sc_hd__mux2_2 _6241_ (.A0(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[3] ),
    .A1(_2468_),
    .S(_3116_),
    .X(_3120_));
 sky130_fd_sc_hd__buf_1 _6242_ (.A(_3120_),
    .X(_0676_));
 sky130_fd_sc_hd__mux2_2 _6243_ (.A0(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[4] ),
    .A1(_2490_),
    .S(_3116_),
    .X(_3121_));
 sky130_fd_sc_hd__buf_1 _6244_ (.A(_3121_),
    .X(_0677_));
 sky130_fd_sc_hd__mux2_2 _6245_ (.A0(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[5] ),
    .A1(_2477_),
    .S(_3116_),
    .X(_3122_));
 sky130_fd_sc_hd__buf_1 _6246_ (.A(_3122_),
    .X(_0678_));
 sky130_fd_sc_hd__mux2_2 _6247_ (.A0(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[6] ),
    .A1(_2474_),
    .S(_3116_),
    .X(_3123_));
 sky130_fd_sc_hd__buf_1 _6248_ (.A(_3123_),
    .X(_0679_));
 sky130_fd_sc_hd__mux2_2 _6249_ (.A0(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[7] ),
    .A1(_2475_),
    .S(_3116_),
    .X(_3124_));
 sky130_fd_sc_hd__buf_1 _6250_ (.A(_3124_),
    .X(_0680_));
 sky130_fd_sc_hd__nor2_2 _6251_ (.A(_2998_),
    .B(_3010_),
    .Y(_0681_));
 sky130_fd_sc_hd__buf_1 _6252_ (.A(_3007_),
    .X(_3125_));
 sky130_fd_sc_hd__mux2_2 _6253_ (.A0(\tree_instances[5].u_tree.u_tree_weight_rom.cached_data[107] ),
    .A1(\tree_instances[5].u_tree.u_tree_weight_rom.gen_tree_5.u_tree_rom.node_data[107] ),
    .S(_3125_),
    .X(_3126_));
 sky130_fd_sc_hd__buf_1 _6254_ (.A(_3126_),
    .X(_0682_));
 sky130_fd_sc_hd__mux2_2 _6255_ (.A0(\tree_instances[6].u_tree.pipeline_frame_id[0][0] ),
    .A1(_1826_),
    .S(_0038_),
    .X(_3127_));
 sky130_fd_sc_hd__buf_1 _6256_ (.A(_3127_),
    .X(_0683_));
 sky130_fd_sc_hd__mux2_2 _6257_ (.A0(\tree_instances[6].u_tree.pipeline_frame_id[0][1] ),
    .A1(_1829_),
    .S(_0038_),
    .X(_3128_));
 sky130_fd_sc_hd__buf_1 _6258_ (.A(_3128_),
    .X(_0684_));
 sky130_fd_sc_hd__mux2_2 _6259_ (.A0(\tree_instances[6].u_tree.pipeline_frame_id[0][2] ),
    .A1(_2595_),
    .S(_0038_),
    .X(_3129_));
 sky130_fd_sc_hd__buf_1 _6260_ (.A(_3129_),
    .X(_0685_));
 sky130_fd_sc_hd__mux2_2 _6261_ (.A0(\tree_instances[6].u_tree.pipeline_frame_id[0][3] ),
    .A1(_1834_),
    .S(_0038_),
    .X(_3130_));
 sky130_fd_sc_hd__buf_1 _6262_ (.A(_3130_),
    .X(_0686_));
 sky130_fd_sc_hd__mux2_2 _6263_ (.A0(\tree_instances[6].u_tree.pipeline_frame_id[0][4] ),
    .A1(\tree_instances[0].u_tree.frame_id_in[4] ),
    .S(_0038_),
    .X(_3131_));
 sky130_fd_sc_hd__buf_1 _6264_ (.A(_3131_),
    .X(_0687_));
 sky130_fd_sc_hd__buf_1 _6265_ (.A(_0933_),
    .X(_3132_));
 sky130_fd_sc_hd__mux2_2 _6266_ (.A0(\tree_instances[5].u_tree.current_node_data[107] ),
    .A1(\tree_instances[5].u_tree.node_data[107] ),
    .S(_3132_),
    .X(_3133_));
 sky130_fd_sc_hd__buf_1 _6267_ (.A(_3133_),
    .X(_0688_));
 sky130_fd_sc_hd__mux2_2 _6268_ (.A0(\tree_instances[6].u_tree.frame_id_out[0] ),
    .A1(\tree_instances[6].u_tree.pipeline_frame_id[0][0] ),
    .S(_0932_),
    .X(_3134_));
 sky130_fd_sc_hd__buf_1 _6269_ (.A(_3134_),
    .X(_0689_));
 sky130_fd_sc_hd__mux2_2 _6270_ (.A0(\tree_instances[6].u_tree.frame_id_out[1] ),
    .A1(\tree_instances[6].u_tree.pipeline_frame_id[0][1] ),
    .S(_0932_),
    .X(_3135_));
 sky130_fd_sc_hd__buf_1 _6271_ (.A(_3135_),
    .X(_0690_));
 sky130_fd_sc_hd__mux2_2 _6272_ (.A0(\tree_instances[6].u_tree.frame_id_out[2] ),
    .A1(\tree_instances[6].u_tree.pipeline_frame_id[0][2] ),
    .S(_0932_),
    .X(_3136_));
 sky130_fd_sc_hd__buf_1 _6273_ (.A(_3136_),
    .X(_0691_));
 sky130_fd_sc_hd__mux2_2 _6274_ (.A0(\tree_instances[6].u_tree.frame_id_out[3] ),
    .A1(\tree_instances[6].u_tree.pipeline_frame_id[0][3] ),
    .S(_0932_),
    .X(_3137_));
 sky130_fd_sc_hd__buf_1 _6275_ (.A(_3137_),
    .X(_0692_));
 sky130_fd_sc_hd__mux2_2 _6276_ (.A0(\tree_instances[6].u_tree.frame_id_out[4] ),
    .A1(\tree_instances[6].u_tree.pipeline_frame_id[0][4] ),
    .S(\tree_instances[6].u_tree.tree_state[3] ),
    .X(_3138_));
 sky130_fd_sc_hd__buf_1 _6277_ (.A(_3138_),
    .X(_0693_));
 sky130_fd_sc_hd__and2_2 _6278_ (.A(_2456_),
    .B(_3102_),
    .X(_3139_));
 sky130_fd_sc_hd__buf_1 _6279_ (.A(_3139_),
    .X(_0694_));
 sky130_fd_sc_hd__and2_2 _6280_ (.A(_2486_),
    .B(_3102_),
    .X(_3140_));
 sky130_fd_sc_hd__buf_1 _6281_ (.A(_3140_),
    .X(_0695_));
 sky130_fd_sc_hd__and2_2 _6282_ (.A(_2481_),
    .B(_3102_),
    .X(_3141_));
 sky130_fd_sc_hd__buf_1 _6283_ (.A(_3141_),
    .X(_0696_));
 sky130_fd_sc_hd__and2_2 _6284_ (.A(_2468_),
    .B(_3102_),
    .X(_3142_));
 sky130_fd_sc_hd__buf_1 _6285_ (.A(_3142_),
    .X(_0697_));
 sky130_fd_sc_hd__and2_2 _6286_ (.A(_2490_),
    .B(_3102_),
    .X(_3143_));
 sky130_fd_sc_hd__buf_1 _6287_ (.A(_3143_),
    .X(_0698_));
 sky130_fd_sc_hd__and2_2 _6288_ (.A(_2477_),
    .B(_3102_),
    .X(_3144_));
 sky130_fd_sc_hd__buf_1 _6289_ (.A(_3144_),
    .X(_0699_));
 sky130_fd_sc_hd__and2_2 _6290_ (.A(_2474_),
    .B(_3102_),
    .X(_3145_));
 sky130_fd_sc_hd__buf_1 _6291_ (.A(_3145_),
    .X(_0700_));
 sky130_fd_sc_hd__and2_2 _6292_ (.A(_2475_),
    .B(_3101_),
    .X(_3146_));
 sky130_fd_sc_hd__buf_1 _6293_ (.A(_3146_),
    .X(_0701_));
 sky130_fd_sc_hd__and2_2 _6294_ (.A(_0945_),
    .B(_3101_),
    .X(_3147_));
 sky130_fd_sc_hd__buf_1 _6295_ (.A(_3147_),
    .X(_0702_));
 sky130_fd_sc_hd__a22o_2 _6296_ (.A1(_0932_),
    .A2(_3081_),
    .B1(_1811_),
    .B2(\tree_instances[6].u_tree.ready_for_next ),
    .X(_0703_));
 sky130_fd_sc_hd__nand2_2 _6297_ (.A(\tree_instances[5].u_tree.pipeline_valid[0] ),
    .B(\tree_instances[5].u_tree.tree_state[0] ),
    .Y(_3148_));
 sky130_fd_sc_hd__o2bb2a_2 _6298_ (.A1_N(_0903_),
    .A2_N(_3148_),
    .B1(_0036_),
    .B2(\tree_instances[5].u_tree.pipeline_valid[0] ),
    .X(_0704_));
 sky130_fd_sc_hd__dfrtp_2 _6299_ (.CLK(clk),
    .D(_0108_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6300_ (.CLK(clk),
    .D(_0109_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6301_ (.CLK(clk),
    .D(_0110_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6302_ (.CLK(clk),
    .D(_0111_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6303_ (.CLK(clk),
    .D(_0112_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6304_ (.CLK(clk),
    .D(_0113_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6305_ (.CLK(clk),
    .D(_0114_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6306_ (.CLK(clk),
    .D(_0115_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6307_ (.CLK(clk),
    .D(_0116_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6308_ (.CLK(clk),
    .D(_0117_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6309_ (.CLK(clk),
    .D(_0118_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6310_ (.CLK(clk),
    .D(_0119_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6311_ (.CLK(clk),
    .D(_0120_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6312_ (.CLK(clk),
    .D(_0121_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6313_ (.CLK(clk),
    .D(_0122_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6314_ (.CLK(clk),
    .D(_0123_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6315_ (.CLK(clk),
    .D(_0124_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6316_ (.CLK(clk),
    .D(_0125_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6317_ (.CLK(clk),
    .D(_0126_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_current_node[0][8] ));
 sky130_fd_sc_hd__dfstp_2 _6318_ (.CLK(clk),
    .D(_0127_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6319_ (.CLK(clk),
    .D(_0105_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6320_ (.CLK(clk),
    .D(_0128_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6321_ (.CLK(clk),
    .D(_0129_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_prediction[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _6322_ (.CLK(clk),
    .D(_0130_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.cache_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6323_ (.CLK(clk),
    .D(_0131_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6324_ (.CLK(clk),
    .D(_0132_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6325_ (.CLK(clk),
    .D(_0133_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6326_ (.CLK(clk),
    .D(_0134_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6327_ (.CLK(clk),
    .D(_0135_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6328_ (.CLK(clk),
    .D(_0136_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6329_ (.CLK(clk),
    .D(_0137_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6330_ (.CLK(clk),
    .D(_0138_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6331_ (.CLK(clk),
    .D(_0139_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6332_ (.CLK(clk),
    .D(_0140_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6333_ (.CLK(clk),
    .D(_0141_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6334_ (.CLK(clk),
    .D(_0142_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6335_ (.CLK(clk),
    .D(_0143_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6336_ (.CLK(clk),
    .D(_0144_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.read_enable ));
 sky130_fd_sc_hd__dfrtp_2 _6337_ (.CLK(clk),
    .D(_0145_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6338_ (.CLK(clk),
    .D(_0146_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6339_ (.CLK(clk),
    .D(_0147_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6340_ (.CLK(clk),
    .D(_0148_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6341_ (.CLK(clk),
    .D(_0149_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6342_ (.CLK(clk),
    .D(_0150_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.prediction_out ));
 sky130_fd_sc_hd__dfstp_2 _6343_ (.CLK(clk),
    .D(_0151_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6344_ (.CLK(clk),
    .D(_0106_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6345_ (.CLK(clk),
    .D(_0152_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6346_ (.CLK(clk),
    .D(_0153_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6347_ (.CLK(clk),
    .D(_0154_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6348_ (.CLK(clk),
    .D(_0155_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6349_ (.CLK(clk),
    .D(_0156_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6350_ (.CLK(clk),
    .D(_0157_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6351_ (.CLK(clk),
    .D(_0158_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6352_ (.CLK(clk),
    .D(_0159_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6353_ (.CLK(clk),
    .D(_0160_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6354_ (.CLK(clk),
    .D(_0161_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.gen_tree_12.u_tree_rom.node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6355_ (.CLK(clk),
    .D(_0162_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6356_ (.CLK(clk),
    .D(_0163_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6357_ (.CLK(clk),
    .D(_0164_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6358_ (.CLK(clk),
    .D(_0165_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6359_ (.CLK(clk),
    .D(_0166_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6360_ (.CLK(clk),
    .D(_0167_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6361_ (.CLK(clk),
    .D(_0168_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6362_ (.CLK(clk),
    .D(_0169_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6363_ (.CLK(clk),
    .D(_0170_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.cached_addr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6364_ (.CLK(clk),
    .D(_0171_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.cached_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6365_ (.CLK(clk),
    .D(_0172_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6366_ (.CLK(clk),
    .D(_0173_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6367_ (.CLK(clk),
    .D(_0174_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6368_ (.CLK(clk),
    .D(_0175_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6369_ (.CLK(clk),
    .D(_0176_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6370_ (.CLK(clk),
    .D(_0177_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.current_node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6371_ (.CLK(clk),
    .D(_0178_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6372_ (.CLK(clk),
    .D(_0179_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6373_ (.CLK(clk),
    .D(_0180_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6374_ (.CLK(clk),
    .D(_0181_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6375_ (.CLK(clk),
    .D(_0182_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6376_ (.CLK(clk),
    .D(_0183_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6377_ (.CLK(clk),
    .D(_0184_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6378_ (.CLK(clk),
    .D(_0185_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6379_ (.CLK(clk),
    .D(_0186_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6380_ (.CLK(clk),
    .D(_0187_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6381_ (.CLK(clk),
    .D(_0188_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6382_ (.CLK(clk),
    .D(_0189_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6383_ (.CLK(clk),
    .D(_0190_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfstp_2 _6384_ (.CLK(clk),
    .D(_0191_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6385_ (.CLK(clk),
    .D(_0107_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6386_ (.CLK(clk),
    .D(_0192_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfstp_2 _6387_ (.CLK(clk),
    .D(_0071_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6388_ (.CLK(clk),
    .D(_0029_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6389_ (.CLK(clk),
    .D(_0030_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6390_ (.CLK(clk),
    .D(_0072_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6391_ (.CLK(clk),
    .D(_0193_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_prediction[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _6392_ (.CLK(clk),
    .D(_0194_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.cache_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6393_ (.CLK(clk),
    .D(_0195_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6394_ (.CLK(clk),
    .D(_0196_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6395_ (.CLK(clk),
    .D(_0197_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6396_ (.CLK(clk),
    .D(_0198_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6397_ (.CLK(clk),
    .D(_0199_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6398_ (.CLK(clk),
    .D(_0200_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6399_ (.CLK(clk),
    .D(_0201_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6400_ (.CLK(clk),
    .D(_0202_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6401_ (.CLK(clk),
    .D(_0203_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6402_ (.CLK(clk),
    .D(_0204_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6403_ (.CLK(clk),
    .D(_0205_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6404_ (.CLK(clk),
    .D(_0206_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6405_ (.CLK(clk),
    .D(_0207_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6406_ (.CLK(clk),
    .D(_0208_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.read_enable ));
 sky130_fd_sc_hd__dfrtp_2 _6407_ (.CLK(clk),
    .D(_0209_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6408_ (.CLK(clk),
    .D(_0210_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6409_ (.CLK(clk),
    .D(_0211_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6410_ (.CLK(clk),
    .D(_0212_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6411_ (.CLK(clk),
    .D(_0213_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6412_ (.CLK(clk),
    .D(_0214_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.prediction_out ));
 sky130_fd_sc_hd__dfstp_2 _6413_ (.CLK(clk),
    .D(_0215_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6414_ (.CLK(clk),
    .D(_0088_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6415_ (.CLK(clk),
    .D(_0216_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfstp_2 _6416_ (.CLK(clk),
    .D(_0063_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6417_ (.CLK(clk),
    .D(_0021_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6418_ (.CLK(clk),
    .D(_0022_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6419_ (.CLK(clk),
    .D(_0064_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6420_ (.CLK(clk),
    .D(_0217_),
    .Q(\tree_instances[10].u_tree.node_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6421_ (.CLK(clk),
    .D(_0218_),
    .Q(\tree_instances[8].u_tree.u_tree_weight_rom.gen_tree_8.u_tree_rom.node_data[12] ));
 sky130_fd_sc_hd__dfstp_2 _6422_ (.CLK(clk),
    .D(_0073_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6423_ (.CLK(clk),
    .D(_0031_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6424_ (.CLK(clk),
    .D(_0032_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6425_ (.CLK(clk),
    .D(_0074_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6426_ (.CLK(clk),
    .D(_0219_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6427_ (.CLK(clk),
    .D(_0220_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6428_ (.CLK(clk),
    .D(_0221_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6429_ (.CLK(clk),
    .D(_0222_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6430_ (.CLK(clk),
    .D(_0223_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6431_ (.CLK(clk),
    .D(_0224_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6432_ (.CLK(clk),
    .D(_0225_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6433_ (.CLK(clk),
    .D(_0226_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.cached_addr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6434_ (.CLK(clk),
    .D(_0227_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.cached_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6435_ (.CLK(clk),
    .D(_0228_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6436_ (.CLK(clk),
    .D(_0229_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6437_ (.CLK(clk),
    .D(_0230_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6438_ (.CLK(clk),
    .D(_0231_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6439_ (.CLK(clk),
    .D(_0232_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6440_ (.CLK(clk),
    .D(_0233_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.current_node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6441_ (.CLK(clk),
    .D(_0234_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6442_ (.CLK(clk),
    .D(_0235_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6443_ (.CLK(clk),
    .D(_0236_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6444_ (.CLK(clk),
    .D(_0237_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6445_ (.CLK(clk),
    .D(_0238_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6446_ (.CLK(clk),
    .D(_0239_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6447_ (.CLK(clk),
    .D(_0240_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6448_ (.CLK(clk),
    .D(_0241_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6449_ (.CLK(clk),
    .D(_0242_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6450_ (.CLK(clk),
    .D(_0243_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6451_ (.CLK(clk),
    .D(_0244_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6452_ (.CLK(clk),
    .D(_0245_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6453_ (.CLK(clk),
    .D(_0246_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfstp_2 _6454_ (.CLK(clk),
    .D(_0247_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6455_ (.CLK(clk),
    .D(_0089_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfxtp_2 _6456_ (.CLK(clk),
    .D(_0248_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.gen_tree_20.u_tree_rom.node_data[12] ));
 sky130_fd_sc_hd__dfstp_2 _6457_ (.CLK(clk),
    .D(_0075_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6458_ (.CLK(clk),
    .D(_0033_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6459_ (.CLK(clk),
    .D(_0034_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6460_ (.CLK(clk),
    .D(_0076_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6461_ (.CLK(clk),
    .D(_0249_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_prediction[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _6462_ (.CLK(clk),
    .D(_0250_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.cache_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6463_ (.CLK(clk),
    .D(_0251_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6464_ (.CLK(clk),
    .D(_0252_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6465_ (.CLK(clk),
    .D(_0253_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6466_ (.CLK(clk),
    .D(_0254_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6467_ (.CLK(clk),
    .D(_0255_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6468_ (.CLK(clk),
    .D(_0256_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6469_ (.CLK(clk),
    .D(_0257_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6470_ (.CLK(clk),
    .D(_0258_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6471_ (.CLK(clk),
    .D(_0259_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6472_ (.CLK(clk),
    .D(_0260_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6473_ (.CLK(clk),
    .D(_0261_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6474_ (.CLK(clk),
    .D(_0262_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6475_ (.CLK(clk),
    .D(_0263_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6476_ (.CLK(clk),
    .D(_0264_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.read_enable ));
 sky130_fd_sc_hd__dfrtp_2 _6477_ (.CLK(clk),
    .D(_0265_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6478_ (.CLK(clk),
    .D(_0266_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6479_ (.CLK(clk),
    .D(_0267_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6480_ (.CLK(clk),
    .D(_0268_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6481_ (.CLK(clk),
    .D(_0269_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6482_ (.CLK(clk),
    .D(_0270_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.prediction_out ));
 sky130_fd_sc_hd__dfstp_2 _6483_ (.CLK(clk),
    .D(_0271_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6484_ (.CLK(clk),
    .D(_0090_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfstp_2 _6485_ (.CLK(clk),
    .D(_0077_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6486_ (.CLK(clk),
    .D(_0035_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6487_ (.CLK(clk),
    .D(_0036_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6488_ (.CLK(clk),
    .D(_0078_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6489_ (.CLK(clk),
    .D(_0272_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_prediction[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _6490_ (.CLK(clk),
    .D(_0273_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.cache_valid ));
 sky130_fd_sc_hd__dfxtp_2 _6491_ (.CLK(clk),
    .D(_0274_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6492_ (.CLK(clk),
    .D(_0275_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6493_ (.CLK(clk),
    .D(_0276_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6494_ (.CLK(clk),
    .D(_0277_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6495_ (.CLK(clk),
    .D(_0278_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6496_ (.CLK(clk),
    .D(_0279_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6497_ (.CLK(clk),
    .D(_0280_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6498_ (.CLK(clk),
    .D(_0281_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.cached_addr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6499_ (.CLK(clk),
    .D(_0282_),
    .Q(\tree_instances[12].u_tree.u_tree_weight_rom.cached_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6500_ (.CLK(clk),
    .D(_0283_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.gen_tree_13.u_tree_rom.node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6501_ (.CLK(clk),
    .D(_0284_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6502_ (.CLK(clk),
    .D(_0285_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6503_ (.CLK(clk),
    .D(_0286_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6504_ (.CLK(clk),
    .D(_0287_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6505_ (.CLK(clk),
    .D(_0288_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6506_ (.CLK(clk),
    .D(_0289_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6507_ (.CLK(clk),
    .D(_0290_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6508_ (.CLK(clk),
    .D(_0291_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6509_ (.CLK(clk),
    .D(_0292_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6510_ (.CLK(clk),
    .D(_0293_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6511_ (.CLK(clk),
    .D(_0294_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6512_ (.CLK(clk),
    .D(_0295_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6513_ (.CLK(clk),
    .D(_0296_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6514_ (.CLK(clk),
    .D(_0297_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.current_node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6515_ (.CLK(clk),
    .D(_0298_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.read_enable ));
 sky130_fd_sc_hd__dfrtp_2 _6516_ (.CLK(clk),
    .D(_0299_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6517_ (.CLK(clk),
    .D(_0300_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6518_ (.CLK(clk),
    .D(_0301_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6519_ (.CLK(clk),
    .D(_0302_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6520_ (.CLK(clk),
    .D(_0303_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6521_ (.CLK(clk),
    .D(_0304_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.prediction_out ));
 sky130_fd_sc_hd__dfstp_2 _6522_ (.CLK(clk),
    .D(_0305_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6523_ (.CLK(clk),
    .D(_0091_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6524_ (.CLK(clk),
    .D(_0306_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfstp_2 _6525_ (.CLK(clk),
    .D(_0061_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6526_ (.CLK(clk),
    .D(_0019_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6527_ (.CLK(clk),
    .D(_0020_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6528_ (.CLK(clk),
    .D(_0062_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfstp_2 _6529_ (.CLK(clk),
    .D(_0079_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6530_ (.CLK(clk),
    .D(_0037_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6531_ (.CLK(clk),
    .D(_0038_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6532_ (.CLK(clk),
    .D(_0080_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6533_ (.CLK(clk),
    .D(_0307_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6534_ (.CLK(clk),
    .D(_0308_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6535_ (.CLK(clk),
    .D(_0309_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6536_ (.CLK(clk),
    .D(_0310_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6537_ (.CLK(clk),
    .D(_0311_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6538_ (.CLK(clk),
    .D(_0312_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6539_ (.CLK(clk),
    .D(_0313_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6540_ (.CLK(clk),
    .D(_0314_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.cached_addr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6541_ (.CLK(clk),
    .D(_0315_),
    .Q(\tree_instances[13].u_tree.u_tree_weight_rom.cached_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6542_ (.CLK(clk),
    .D(_0316_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6543_ (.CLK(clk),
    .D(_0317_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6544_ (.CLK(clk),
    .D(_0318_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6545_ (.CLK(clk),
    .D(_0319_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6546_ (.CLK(clk),
    .D(_0320_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6547_ (.CLK(clk),
    .D(_0321_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.current_node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6548_ (.CLK(clk),
    .D(_0322_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6549_ (.CLK(clk),
    .D(_0323_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6550_ (.CLK(clk),
    .D(_0324_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6551_ (.CLK(clk),
    .D(_0325_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6552_ (.CLK(clk),
    .D(_0326_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6553_ (.CLK(clk),
    .D(_0327_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6554_ (.CLK(clk),
    .D(_0328_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6555_ (.CLK(clk),
    .D(_0329_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6556_ (.CLK(clk),
    .D(_0330_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6557_ (.CLK(clk),
    .D(_0331_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6558_ (.CLK(clk),
    .D(_0332_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6559_ (.CLK(clk),
    .D(_0333_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6560_ (.CLK(clk),
    .D(_0334_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfstp_2 _6561_ (.CLK(clk),
    .D(_0335_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6562_ (.CLK(clk),
    .D(_0092_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfstp_2 _6563_ (.CLK(clk),
    .D(_0081_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6564_ (.CLK(clk),
    .D(_0039_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6565_ (.CLK(clk),
    .D(_0040_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6566_ (.CLK(clk),
    .D(_0082_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6567_ (.CLK(clk),
    .D(_0336_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6568_ (.CLK(clk),
    .D(_0337_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6569_ (.CLK(clk),
    .D(_0338_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6570_ (.CLK(clk),
    .D(_0339_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6571_ (.CLK(clk),
    .D(_0340_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6572_ (.CLK(clk),
    .D(_0341_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6573_ (.CLK(clk),
    .D(_0342_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6574_ (.CLK(clk),
    .D(_0343_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6575_ (.CLK(clk),
    .D(_0344_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6576_ (.CLK(clk),
    .D(_0345_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6577_ (.CLK(clk),
    .D(_0346_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6578_ (.CLK(clk),
    .D(_0347_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6579_ (.CLK(clk),
    .D(_0348_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6580_ (.CLK(clk),
    .D(_0349_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6581_ (.CLK(clk),
    .D(_0350_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6582_ (.CLK(clk),
    .D(_0351_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6583_ (.CLK(clk),
    .D(_0352_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6584_ (.CLK(clk),
    .D(_0353_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfstp_2 _6585_ (.CLK(clk),
    .D(_0354_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6586_ (.CLK(clk),
    .D(_0093_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfstp_2 _6587_ (.CLK(clk),
    .D(_0083_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6588_ (.CLK(clk),
    .D(_0041_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6589_ (.CLK(clk),
    .D(_0042_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6590_ (.CLK(clk),
    .D(_0084_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6591_ (.CLK(clk),
    .D(_0355_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_prediction[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _6592_ (.CLK(clk),
    .D(_0356_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.cache_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6593_ (.CLK(clk),
    .D(_0357_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6594_ (.CLK(clk),
    .D(_0358_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6595_ (.CLK(clk),
    .D(_0359_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6596_ (.CLK(clk),
    .D(_0360_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6597_ (.CLK(clk),
    .D(_0361_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6598_ (.CLK(clk),
    .D(_0362_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6599_ (.CLK(clk),
    .D(_0363_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6600_ (.CLK(clk),
    .D(_0364_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6601_ (.CLK(clk),
    .D(_0365_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6602_ (.CLK(clk),
    .D(_0366_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6603_ (.CLK(clk),
    .D(_0367_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6604_ (.CLK(clk),
    .D(_0368_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6605_ (.CLK(clk),
    .D(_0369_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6606_ (.CLK(clk),
    .D(_0370_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.read_enable ));
 sky130_fd_sc_hd__dfrtp_2 _6607_ (.CLK(clk),
    .D(_0371_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6608_ (.CLK(clk),
    .D(_0372_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6609_ (.CLK(clk),
    .D(_0373_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6610_ (.CLK(clk),
    .D(_0374_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6611_ (.CLK(clk),
    .D(_0375_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6612_ (.CLK(clk),
    .D(_0376_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.prediction_out ));
 sky130_fd_sc_hd__dfstp_2 _6613_ (.CLK(clk),
    .D(_0377_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6614_ (.CLK(clk),
    .D(_0094_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6615_ (.CLK(clk),
    .D(_0378_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6616_ (.CLK(clk),
    .D(_0379_),
    .Q(\tree_instances[10].u_tree.u_tree_weight_rom.gen_tree_10.u_tree_rom.node_data[12] ));
 sky130_fd_sc_hd__dfstp_2 _6617_ (.CLK(clk),
    .D(_0085_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6618_ (.CLK(clk),
    .D(_0043_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6619_ (.CLK(clk),
    .D(_0044_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6620_ (.CLK(clk),
    .D(_0086_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6621_ (.CLK(clk),
    .D(_0380_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.cached_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6622_ (.CLK(clk),
    .D(_0381_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6623_ (.CLK(clk),
    .D(_0382_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6624_ (.CLK(clk),
    .D(_0383_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6625_ (.CLK(clk),
    .D(_0384_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6626_ (.CLK(clk),
    .D(_0385_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6627_ (.CLK(clk),
    .D(_0386_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6628_ (.CLK(clk),
    .D(_0387_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6629_ (.CLK(clk),
    .D(_0388_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6630_ (.CLK(clk),
    .D(_0389_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_current_node[0][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6631_ (.CLK(clk),
    .D(_0390_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6632_ (.CLK(clk),
    .D(_0391_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6633_ (.CLK(clk),
    .D(_0392_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6634_ (.CLK(clk),
    .D(_0393_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6635_ (.CLK(clk),
    .D(_0394_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6636_ (.CLK(clk),
    .D(_0395_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.current_node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6637_ (.CLK(clk),
    .D(_0396_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6638_ (.CLK(clk),
    .D(_0397_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6639_ (.CLK(clk),
    .D(_0398_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6640_ (.CLK(clk),
    .D(_0399_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6641_ (.CLK(clk),
    .D(_0400_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6642_ (.CLK(clk),
    .D(_0401_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6643_ (.CLK(clk),
    .D(_0402_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6644_ (.CLK(clk),
    .D(_0403_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6645_ (.CLK(clk),
    .D(_0404_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6646_ (.CLK(clk),
    .D(_0405_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6647_ (.CLK(clk),
    .D(_0406_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6648_ (.CLK(clk),
    .D(_0407_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6649_ (.CLK(clk),
    .D(_0408_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfstp_2 _6650_ (.CLK(clk),
    .D(_0409_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6651_ (.CLK(clk),
    .D(_0095_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfstp_2 _6652_ (.CLK(clk),
    .D(_0059_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6653_ (.CLK(clk),
    .D(_0017_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6654_ (.CLK(clk),
    .D(_0018_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6655_ (.CLK(clk),
    .D(_0060_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6656_ (.CLK(clk),
    .D(_0410_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[9].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfstp_2 _6657_ (.CLK(clk),
    .D(_0053_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6658_ (.CLK(clk),
    .D(_0011_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6659_ (.CLK(clk),
    .D(_0012_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6660_ (.CLK(clk),
    .D(_0054_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[13].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6661_ (.CLK(clk),
    .D(_0411_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6662_ (.CLK(clk),
    .D(_0412_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6663_ (.CLK(clk),
    .D(_0413_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6664_ (.CLK(clk),
    .D(_0414_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6665_ (.CLK(clk),
    .D(_0415_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6666_ (.CLK(clk),
    .D(_0416_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6667_ (.CLK(clk),
    .D(_0417_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6668_ (.CLK(clk),
    .D(_0418_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.cached_addr[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6669_ (.CLK(clk),
    .D(_0419_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6670_ (.CLK(clk),
    .D(_0420_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6671_ (.CLK(clk),
    .D(_0421_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6672_ (.CLK(clk),
    .D(_0422_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6673_ (.CLK(clk),
    .D(_0423_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6674_ (.CLK(clk),
    .D(_0424_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6675_ (.CLK(clk),
    .D(_0425_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6676_ (.CLK(clk),
    .D(_0426_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6677_ (.CLK(clk),
    .D(_0427_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6678_ (.CLK(clk),
    .D(_0428_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfstp_2 _6679_ (.CLK(clk),
    .D(_0429_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6680_ (.CLK(clk),
    .D(_0096_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6681_ (.CLK(clk),
    .D(_0430_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6682_ (.CLK(clk),
    .D(_0431_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6683_ (.CLK(clk),
    .D(_0432_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6684_ (.CLK(clk),
    .D(_0433_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6685_ (.CLK(clk),
    .D(_0434_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6686_ (.CLK(clk),
    .D(_0435_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6687_ (.CLK(clk),
    .D(_0436_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6688_ (.CLK(clk),
    .D(_0437_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6689_ (.CLK(clk),
    .D(_0438_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6690_ (.CLK(clk),
    .D(_0439_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6691_ (.CLK(clk),
    .D(_0440_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6692_ (.CLK(clk),
    .D(_0441_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6693_ (.CLK(clk),
    .D(_0442_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6694_ (.CLK(clk),
    .D(_0443_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6695_ (.CLK(clk),
    .D(_0444_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6696_ (.CLK(clk),
    .D(_0445_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6697_ (.CLK(clk),
    .D(_0446_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6698_ (.CLK(clk),
    .D(_0447_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6699_ (.CLK(clk),
    .D(_0448_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[18].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfstp_2 _6700_ (.CLK(clk),
    .D(_0449_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6701_ (.CLK(clk),
    .D(_0097_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6702_ (.CLK(clk),
    .D(_0450_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6703_ (.CLK(clk),
    .D(_0451_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6704_ (.CLK(clk),
    .D(_0452_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[8].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6705_ (.CLK(clk),
    .D(_0453_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6706_ (.CLK(clk),
    .D(_0454_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6707_ (.CLK(clk),
    .D(_0455_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_prediction[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _6708_ (.CLK(clk),
    .D(_0456_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.cache_valid ));
 sky130_fd_sc_hd__dfxtp_2 _6709_ (.CLK(clk),
    .D(_0457_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6710_ (.CLK(clk),
    .D(_0458_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6711_ (.CLK(clk),
    .D(_0459_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6712_ (.CLK(clk),
    .D(_0460_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6713_ (.CLK(clk),
    .D(_0461_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6714_ (.CLK(clk),
    .D(_0462_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6715_ (.CLK(clk),
    .D(_0463_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6716_ (.CLK(clk),
    .D(_0464_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.cached_addr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6717_ (.CLK(clk),
    .D(_0465_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.cached_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6718_ (.CLK(clk),
    .D(_0466_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6719_ (.CLK(clk),
    .D(_0467_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6720_ (.CLK(clk),
    .D(_0468_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6721_ (.CLK(clk),
    .D(_0469_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6722_ (.CLK(clk),
    .D(_0470_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6723_ (.CLK(clk),
    .D(_0471_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6724_ (.CLK(clk),
    .D(_0472_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6725_ (.CLK(clk),
    .D(_0473_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6726_ (.CLK(clk),
    .D(_0474_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6727_ (.CLK(clk),
    .D(_0475_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6728_ (.CLK(clk),
    .D(_0476_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6729_ (.CLK(clk),
    .D(_0477_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6730_ (.CLK(clk),
    .D(_0478_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6731_ (.CLK(clk),
    .D(_0479_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.current_node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6732_ (.CLK(clk),
    .D(_0480_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.read_enable ));
 sky130_fd_sc_hd__dfrtp_2 _6733_ (.CLK(clk),
    .D(_0481_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6734_ (.CLK(clk),
    .D(_0482_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6735_ (.CLK(clk),
    .D(_0483_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6736_ (.CLK(clk),
    .D(_0484_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6737_ (.CLK(clk),
    .D(_0485_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6738_ (.CLK(clk),
    .D(_0486_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.prediction_out ));
 sky130_fd_sc_hd__dfstp_2 _6739_ (.CLK(clk),
    .D(_0487_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6740_ (.CLK(clk),
    .D(_0099_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6741_ (.CLK(clk),
    .D(_0488_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[16].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfstp_2 _6742_ (.CLK(clk),
    .D(_0057_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6743_ (.CLK(clk),
    .D(_0015_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6744_ (.CLK(clk),
    .D(_0016_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6745_ (.CLK(clk),
    .D(_0058_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[15].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6746_ (.CLK(clk),
    .D(_0489_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.gen_tree_3.u_tree_rom.node_data[107] ));
 sky130_fd_sc_hd__dfxtp_2 _6747_ (.CLK(clk),
    .D(_0490_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.gen_tree_5.u_tree_rom.node_data[107] ));
 sky130_fd_sc_hd__dfstp_2 _6748_ (.CLK(clk),
    .D(_0047_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6749_ (.CLK(clk),
    .D(_0005_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6750_ (.CLK(clk),
    .D(_0006_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6751_ (.CLK(clk),
    .D(_0048_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[10].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfstp_2 _6752_ (.CLK(clk),
    .D(_0049_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6753_ (.CLK(clk),
    .D(_0007_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6754_ (.CLK(clk),
    .D(_0008_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6755_ (.CLK(clk),
    .D(_0050_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6756_ (.CLK(clk),
    .D(_0491_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[11].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6757_ (.CLK(clk),
    .D(_0492_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6758_ (.CLK(clk),
    .D(_0493_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6759_ (.CLK(clk),
    .D(_0000_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(prediction_valid));
 sky130_fd_sc_hd__dfrtp_2 _6760_ (.CLK(clk),
    .D(_0494_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(prediction_out));
 sky130_fd_sc_hd__dfrtp_2 _6761_ (.CLK(clk),
    .D(_0495_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(frame_id_out[0]));
 sky130_fd_sc_hd__dfrtp_2 _6762_ (.CLK(clk),
    .D(_0496_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(frame_id_out[1]));
 sky130_fd_sc_hd__dfrtp_2 _6763_ (.CLK(clk),
    .D(_0497_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(frame_id_out[2]));
 sky130_fd_sc_hd__dfrtp_2 _6764_ (.CLK(clk),
    .D(_0498_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(frame_id_out[3]));
 sky130_fd_sc_hd__dfrtp_2 _6765_ (.CLK(clk),
    .D(_0499_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(frame_id_out[4]));
 sky130_fd_sc_hd__dfrtp_2 _6766_ (.CLK(clk),
    .D(_0500_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.frame_id_in[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6767_ (.CLK(clk),
    .D(_0501_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.frame_id_in[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6768_ (.CLK(clk),
    .D(_0502_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.frame_id_in[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6769_ (.CLK(clk),
    .D(_0503_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.frame_id_in[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6770_ (.CLK(clk),
    .D(_0504_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.frame_id_in[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6771_ (.CLK(clk),
    .D(_0505_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\attack_votes[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6772_ (.CLK(clk),
    .D(_0506_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\attack_votes[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6773_ (.CLK(clk),
    .D(_0507_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\attack_votes[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6774_ (.CLK(clk),
    .D(_0508_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\attack_votes[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6775_ (.CLK(clk),
    .D(_0509_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\attack_votes[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6776_ (.CLK(clk),
    .D(_0510_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\complete_votes[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6777_ (.CLK(clk),
    .D(_0511_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\complete_votes[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6778_ (.CLK(clk),
    .D(_0512_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\complete_votes[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6779_ (.CLK(clk),
    .D(_0513_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\complete_votes[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6780_ (.CLK(clk),
    .D(_0514_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\complete_votes[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6781_ (.CLK(clk),
    .D(_0515_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\current_voting_frame[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6782_ (.CLK(clk),
    .D(_0516_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\current_voting_frame[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6783_ (.CLK(clk),
    .D(_0517_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\current_voting_frame[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6784_ (.CLK(clk),
    .D(_0518_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\current_voting_frame[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6785_ (.CLK(clk),
    .D(_0519_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\current_voting_frame[4] ));
 sky130_fd_sc_hd__dfstp_2 _6786_ (.CLK(clk),
    .D(_0069_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6787_ (.CLK(clk),
    .D(_0027_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6788_ (.CLK(clk),
    .D(_0028_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6789_ (.CLK(clk),
    .D(_0070_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfstp_2 _6790_ (.CLK(clk),
    .D(_0045_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6791_ (.CLK(clk),
    .D(_0003_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6792_ (.CLK(clk),
    .D(_0004_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6793_ (.CLK(clk),
    .D(_0046_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfstp_2 _6794_ (.CLK(clk),
    .D(_0051_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6795_ (.CLK(clk),
    .D(_0009_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6796_ (.CLK(clk),
    .D(_0010_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6797_ (.CLK(clk),
    .D(_0052_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[12].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6798_ (.CLK(clk),
    .D(_0520_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6799_ (.CLK(clk),
    .D(_0521_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6800_ (.CLK(clk),
    .D(_0522_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6801_ (.CLK(clk),
    .D(_0523_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6802_ (.CLK(clk),
    .D(_0524_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6803_ (.CLK(clk),
    .D(_0525_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6804_ (.CLK(clk),
    .D(_0526_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6805_ (.CLK(clk),
    .D(_0527_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6806_ (.CLK(clk),
    .D(_0528_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6807_ (.CLK(clk),
    .D(_0529_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfstp_2 _6808_ (.CLK(clk),
    .D(_0530_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6809_ (.CLK(clk),
    .D(_0087_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[0].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfxtp_2 _6810_ (.CLK(clk),
    .D(_0531_),
    .Q(\tree_instances[8].u_tree.node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6811_ (.CLK(clk),
    .D(_0532_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_prediction[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _6812_ (.CLK(clk),
    .D(_0533_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.cache_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6813_ (.CLK(clk),
    .D(_0534_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6814_ (.CLK(clk),
    .D(_0535_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6815_ (.CLK(clk),
    .D(_0536_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6816_ (.CLK(clk),
    .D(_0537_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6817_ (.CLK(clk),
    .D(_0538_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6818_ (.CLK(clk),
    .D(_0539_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6819_ (.CLK(clk),
    .D(_0540_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6820_ (.CLK(clk),
    .D(_0541_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6821_ (.CLK(clk),
    .D(_0542_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6822_ (.CLK(clk),
    .D(_0543_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6823_ (.CLK(clk),
    .D(_0544_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6824_ (.CLK(clk),
    .D(_0545_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6825_ (.CLK(clk),
    .D(_0546_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6826_ (.CLK(clk),
    .D(_0547_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.read_enable ));
 sky130_fd_sc_hd__dfrtp_2 _6827_ (.CLK(clk),
    .D(_0548_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6828_ (.CLK(clk),
    .D(_0549_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6829_ (.CLK(clk),
    .D(_0550_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6830_ (.CLK(clk),
    .D(_0551_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6831_ (.CLK(clk),
    .D(_0552_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6832_ (.CLK(clk),
    .D(_0553_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.prediction_out ));
 sky130_fd_sc_hd__dfstp_2 _6833_ (.CLK(clk),
    .D(_0554_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6834_ (.CLK(clk),
    .D(_0098_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfxtp_2 _6835_ (.CLK(clk),
    .D(_0555_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.cached_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6836_ (.CLK(clk),
    .D(_0556_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6837_ (.CLK(clk),
    .D(_0557_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6838_ (.CLK(clk),
    .D(_0558_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6839_ (.CLK(clk),
    .D(_0559_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6840_ (.CLK(clk),
    .D(_0560_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6841_ (.CLK(clk),
    .D(_0561_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6842_ (.CLK(clk),
    .D(_0562_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6843_ (.CLK(clk),
    .D(_0563_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6844_ (.CLK(clk),
    .D(_0564_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_current_node[0][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6845_ (.CLK(clk),
    .D(_0565_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_current_node[0][9] ));
 sky130_fd_sc_hd__dfrtp_2 _6846_ (.CLK(clk),
    .D(_0566_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6847_ (.CLK(clk),
    .D(_0567_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6848_ (.CLK(clk),
    .D(_0568_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6849_ (.CLK(clk),
    .D(_0569_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6850_ (.CLK(clk),
    .D(_0570_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6851_ (.CLK(clk),
    .D(_0571_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.current_node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6852_ (.CLK(clk),
    .D(_0572_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6853_ (.CLK(clk),
    .D(_0573_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6854_ (.CLK(clk),
    .D(_0574_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6855_ (.CLK(clk),
    .D(_0575_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6856_ (.CLK(clk),
    .D(_0576_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6857_ (.CLK(clk),
    .D(_0577_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6858_ (.CLK(clk),
    .D(_0578_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6859_ (.CLK(clk),
    .D(_0579_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6860_ (.CLK(clk),
    .D(_0580_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6861_ (.CLK(clk),
    .D(_0581_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6862_ (.CLK(clk),
    .D(_0582_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6863_ (.CLK(clk),
    .D(_0583_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6864_ (.CLK(clk),
    .D(_0584_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[20].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfstp_2 _6865_ (.CLK(clk),
    .D(_0585_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6866_ (.CLK(clk),
    .D(_0100_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[2].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6867_ (.CLK(clk),
    .D(_0586_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[7].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6868_ (.CLK(clk),
    .D(_0587_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_prediction[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _6869_ (.CLK(clk),
    .D(_0588_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.cache_valid ));
 sky130_fd_sc_hd__dfxtp_2 _6870_ (.CLK(clk),
    .D(_0589_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6871_ (.CLK(clk),
    .D(_0590_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6872_ (.CLK(clk),
    .D(_0591_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6873_ (.CLK(clk),
    .D(_0592_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6874_ (.CLK(clk),
    .D(_0593_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6875_ (.CLK(clk),
    .D(_0594_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6876_ (.CLK(clk),
    .D(_0595_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6877_ (.CLK(clk),
    .D(_0596_),
    .Q(\tree_instances[20].u_tree.u_tree_weight_rom.cached_addr[7] ));
 sky130_fd_sc_hd__dfrtp_2 _6878_ (.CLK(clk),
    .D(_0597_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6879_ (.CLK(clk),
    .D(_0598_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6880_ (.CLK(clk),
    .D(_0599_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6881_ (.CLK(clk),
    .D(_0600_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6882_ (.CLK(clk),
    .D(_0601_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6883_ (.CLK(clk),
    .D(_0602_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.read_enable ));
 sky130_fd_sc_hd__dfrtp_2 _6884_ (.CLK(clk),
    .D(_0603_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6885_ (.CLK(clk),
    .D(_0604_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6886_ (.CLK(clk),
    .D(_0605_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6887_ (.CLK(clk),
    .D(_0606_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6888_ (.CLK(clk),
    .D(_0607_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6889_ (.CLK(clk),
    .D(_0608_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.prediction_out ));
 sky130_fd_sc_hd__dfstp_2 _6890_ (.CLK(clk),
    .D(_0609_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6891_ (.CLK(clk),
    .D(_0101_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfstp_2 _6892_ (.CLK(clk),
    .D(_0067_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6893_ (.CLK(clk),
    .D(_0025_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6894_ (.CLK(clk),
    .D(_0026_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6895_ (.CLK(clk),
    .D(_0068_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6896_ (.CLK(clk),
    .D(_0610_),
    .Q(\tree_instances[1].u_tree.node_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6897_ (.CLK(clk),
    .D(_0611_),
    .Q(\tree_instances[3].u_tree.node_data[107] ));
 sky130_fd_sc_hd__dfxtp_2 _6898_ (.CLK(clk),
    .D(_0612_),
    .Q(\tree_instances[5].u_tree.node_data[107] ));
 sky130_fd_sc_hd__dfxtp_2 _6899_ (.CLK(clk),
    .D(_0001_),
    .Q(\tree_instances[16].u_tree.u_tree_weight_rom.gen_tree_16.u_tree_rom.node_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6900_ (.CLK(clk),
    .D(_0613_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6901_ (.CLK(clk),
    .D(_0614_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6902_ (.CLK(clk),
    .D(_0615_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6903_ (.CLK(clk),
    .D(_0616_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6904_ (.CLK(clk),
    .D(_0617_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6905_ (.CLK(clk),
    .D(_0618_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6906_ (.CLK(clk),
    .D(_0619_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6907_ (.CLK(clk),
    .D(_0620_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.cached_addr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6908_ (.CLK(clk),
    .D(_0621_),
    .Q(\tree_instances[3].u_tree.u_tree_weight_rom.cached_data[107] ));
 sky130_fd_sc_hd__dfrtp_2 _6909_ (.CLK(clk),
    .D(_0622_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6910_ (.CLK(clk),
    .D(_0623_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6911_ (.CLK(clk),
    .D(_0624_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6912_ (.CLK(clk),
    .D(_0625_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6913_ (.CLK(clk),
    .D(_0626_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6914_ (.CLK(clk),
    .D(_0627_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.current_node_data[107] ));
 sky130_fd_sc_hd__dfrtp_2 _6915_ (.CLK(clk),
    .D(_0628_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6916_ (.CLK(clk),
    .D(_0629_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6917_ (.CLK(clk),
    .D(_0630_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6918_ (.CLK(clk),
    .D(_0631_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6919_ (.CLK(clk),
    .D(_0632_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6920_ (.CLK(clk),
    .D(_0633_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6921_ (.CLK(clk),
    .D(_0634_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6922_ (.CLK(clk),
    .D(_0635_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6923_ (.CLK(clk),
    .D(_0636_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6924_ (.CLK(clk),
    .D(_0637_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6925_ (.CLK(clk),
    .D(_0638_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6926_ (.CLK(clk),
    .D(_0639_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6927_ (.CLK(clk),
    .D(_0640_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[3].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfstp_2 _6928_ (.CLK(clk),
    .D(_0641_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6929_ (.CLK(clk),
    .D(_0102_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6930_ (.CLK(clk),
    .D(_0642_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[17].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6931_ (.CLK(clk),
    .D(_0643_),
    .Q(\tree_instances[12].u_tree.node_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6932_ (.CLK(clk),
    .D(_0644_),
    .Q(\tree_instances[13].u_tree.node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6933_ (.CLK(clk),
    .D(_0645_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[1].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6934_ (.CLK(clk),
    .D(_0646_),
    .Q(\tree_instances[20].u_tree.node_data[12] ));
 sky130_fd_sc_hd__dfrtp_2 _6935_ (.CLK(clk),
    .D(_0647_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6936_ (.CLK(clk),
    .D(_0648_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_prediction[0][0] ));
 sky130_fd_sc_hd__dfxtp_2 _6937_ (.CLK(clk),
    .D(_0649_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cache_valid ));
 sky130_fd_sc_hd__dfrtp_2 _6938_ (.CLK(clk),
    .D(_0650_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6939_ (.CLK(clk),
    .D(_0651_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6940_ (.CLK(clk),
    .D(_0652_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6941_ (.CLK(clk),
    .D(_0653_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6942_ (.CLK(clk),
    .D(_0654_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6943_ (.CLK(clk),
    .D(_0655_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6944_ (.CLK(clk),
    .D(_0656_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6945_ (.CLK(clk),
    .D(_0657_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6946_ (.CLK(clk),
    .D(_0658_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[4].u_tree.pipeline_current_node[0][8] ));
 sky130_fd_sc_hd__dfrtp_2 _6947_ (.CLK(clk),
    .D(_0659_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6948_ (.CLK(clk),
    .D(_0660_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6949_ (.CLK(clk),
    .D(_0661_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6950_ (.CLK(clk),
    .D(_0662_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6951_ (.CLK(clk),
    .D(_0663_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6952_ (.CLK(clk),
    .D(_0664_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.read_enable ));
 sky130_fd_sc_hd__dfrtp_2 _6953_ (.CLK(clk),
    .D(_0665_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6954_ (.CLK(clk),
    .D(_0666_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6955_ (.CLK(clk),
    .D(_0667_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6956_ (.CLK(clk),
    .D(_0668_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6957_ (.CLK(clk),
    .D(_0669_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6958_ (.CLK(clk),
    .D(_0670_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.prediction_out ));
 sky130_fd_sc_hd__dfstp_2 _6959_ (.CLK(clk),
    .D(_0671_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6960_ (.CLK(clk),
    .D(_0103_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfxtp_2 _6961_ (.CLK(clk),
    .D(_0672_),
    .Q(\tree_instances[16].u_tree.node_data[12] ));
 sky130_fd_sc_hd__dfstp_2 _6962_ (.CLK(clk),
    .D(_0055_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6963_ (.CLK(clk),
    .D(_0013_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6964_ (.CLK(clk),
    .D(_0014_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6965_ (.CLK(clk),
    .D(_0056_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[14].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6966_ (.CLK(clk),
    .D(_0002_),
    .Q(\tree_instances[1].u_tree.u_tree_weight_rom.gen_tree_1.u_tree_rom.node_data[12] ));
 sky130_fd_sc_hd__dfxtp_2 _6967_ (.CLK(clk),
    .D(_0673_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[0] ));
 sky130_fd_sc_hd__dfxtp_2 _6968_ (.CLK(clk),
    .D(_0674_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[1] ));
 sky130_fd_sc_hd__dfxtp_2 _6969_ (.CLK(clk),
    .D(_0675_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[2] ));
 sky130_fd_sc_hd__dfxtp_2 _6970_ (.CLK(clk),
    .D(_0676_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[3] ));
 sky130_fd_sc_hd__dfxtp_2 _6971_ (.CLK(clk),
    .D(_0677_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[4] ));
 sky130_fd_sc_hd__dfxtp_2 _6972_ (.CLK(clk),
    .D(_0678_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[5] ));
 sky130_fd_sc_hd__dfxtp_2 _6973_ (.CLK(clk),
    .D(_0679_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[6] ));
 sky130_fd_sc_hd__dfxtp_2 _6974_ (.CLK(clk),
    .D(_0680_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[7] ));
 sky130_fd_sc_hd__dfxtp_2 _6975_ (.CLK(clk),
    .D(_0681_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cached_addr[8] ));
 sky130_fd_sc_hd__dfxtp_2 _6976_ (.CLK(clk),
    .D(_0682_),
    .Q(\tree_instances[5].u_tree.u_tree_weight_rom.cached_data[107] ));
 sky130_fd_sc_hd__dfrtp_2 _6977_ (.CLK(clk),
    .D(_0683_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_frame_id[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6978_ (.CLK(clk),
    .D(_0684_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_frame_id[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6979_ (.CLK(clk),
    .D(_0685_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_frame_id[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6980_ (.CLK(clk),
    .D(_0686_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_frame_id[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6981_ (.CLK(clk),
    .D(_0687_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.pipeline_frame_id[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6982_ (.CLK(clk),
    .D(_0688_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.current_node_data[107] ));
 sky130_fd_sc_hd__dfrtp_2 _6983_ (.CLK(clk),
    .D(_0689_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.frame_id_out[0] ));
 sky130_fd_sc_hd__dfrtp_2 _6984_ (.CLK(clk),
    .D(_0690_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.frame_id_out[1] ));
 sky130_fd_sc_hd__dfrtp_2 _6985_ (.CLK(clk),
    .D(_0691_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.frame_id_out[2] ));
 sky130_fd_sc_hd__dfrtp_2 _6986_ (.CLK(clk),
    .D(_0692_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.frame_id_out[3] ));
 sky130_fd_sc_hd__dfrtp_2 _6987_ (.CLK(clk),
    .D(_0693_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.frame_id_out[4] ));
 sky130_fd_sc_hd__dfrtp_2 _6988_ (.CLK(clk),
    .D(_0694_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_current_node[0][0] ));
 sky130_fd_sc_hd__dfrtp_2 _6989_ (.CLK(clk),
    .D(_0695_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_current_node[0][1] ));
 sky130_fd_sc_hd__dfrtp_2 _6990_ (.CLK(clk),
    .D(_0696_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_current_node[0][2] ));
 sky130_fd_sc_hd__dfrtp_2 _6991_ (.CLK(clk),
    .D(_0697_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_current_node[0][3] ));
 sky130_fd_sc_hd__dfrtp_2 _6992_ (.CLK(clk),
    .D(_0698_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_current_node[0][4] ));
 sky130_fd_sc_hd__dfrtp_2 _6993_ (.CLK(clk),
    .D(_0699_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_current_node[0][5] ));
 sky130_fd_sc_hd__dfrtp_2 _6994_ (.CLK(clk),
    .D(_0700_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_current_node[0][6] ));
 sky130_fd_sc_hd__dfrtp_2 _6995_ (.CLK(clk),
    .D(_0701_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_current_node[0][7] ));
 sky130_fd_sc_hd__dfrtp_2 _6996_ (.CLK(clk),
    .D(_0702_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_current_node[0][8] ));
 sky130_fd_sc_hd__dfstp_2 _6997_ (.CLK(clk),
    .D(_0703_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.ready_for_next ));
 sky130_fd_sc_hd__dfrtp_2 _6998_ (.CLK(clk),
    .D(_0104_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[6].u_tree.prediction_valid ));
 sky130_fd_sc_hd__dfstp_2 _6999_ (.CLK(clk),
    .D(_0065_),
    .SET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.tree_state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7000_ (.CLK(clk),
    .D(_0023_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.tree_state[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7001_ (.CLK(clk),
    .D(_0024_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.tree_state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7002_ (.CLK(clk),
    .D(_0066_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[19].u_tree.tree_state[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7003_ (.CLK(clk),
    .D(_0704_),
    .RESET_B(\tree_instances[0].u_tree.rst_n ),
    .Q(\tree_instances[5].u_tree.pipeline_valid[0] ));
 sky130_fd_sc_hd__clkbuf_16 rst_buf (.A(rst_n),
    .X(\tree_instances[0].u_tree.rst_n ));
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Right_0 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Right_1 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Right_2 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Right_3 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Right_4 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Right_5 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Right_6 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Right_7 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Right_8 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Right_9 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Right_10 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Right_11 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Right_12 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Right_13 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Right_14 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Right_15 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Right_16 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Right_17 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Right_18 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Right_19 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Right_20 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Right_21 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Right_22 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Right_23 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Right_24 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Right_25 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Right_26 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Right_27 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Right_28 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Right_29 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Right_30 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Right_31 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Right_32 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Right_33 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Right_34 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Right_35 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Right_36 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Right_37 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Right_38 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Right_39 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Right_40 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Right_41 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Right_42 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Right_43 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Right_44 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Right_45 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Right_46 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Right_47 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Right_48 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Right_49 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Right_50 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Right_51 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Right_52 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Right_53 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Right_54 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Right_55 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Right_56 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Right_57 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Right_58 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Right_59 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Right_60 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Right_61 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Right_62 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Right_63 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Right_64 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Right_65 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Right_66 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Right_67 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Right_68 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Right_69 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Right_70 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Right_71 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Right_72 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Right_73 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Right_74 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Right_75 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Right_76 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Right_77 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Right_78 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Right_79 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Right_80 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Right_81 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Right_82 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Right_83 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Right_84 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Right_85 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Right_86 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Right_87 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Right_88 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Right_89 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Right_90 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Right_91 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Right_92 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Right_93 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Right_94 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Right_95 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Right_96 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Right_97 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Right_98 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Right_99 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Right_100 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Right_101 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Right_102 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Right_103 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Right_104 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Right_105 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Right_106 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Right_107 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Right_108 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Right_109 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Right_110 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Right_111 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_0_Left_112 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_1_Left_113 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_2_Left_114 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_3_Left_115 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_4_Left_116 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_5_Left_117 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_6_Left_118 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_7_Left_119 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_8_Left_120 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_9_Left_121 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_10_Left_122 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_11_Left_123 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_12_Left_124 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_13_Left_125 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_14_Left_126 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_15_Left_127 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_16_Left_128 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_17_Left_129 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_18_Left_130 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_19_Left_131 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_20_Left_132 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_21_Left_133 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_22_Left_134 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_23_Left_135 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_24_Left_136 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_25_Left_137 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_26_Left_138 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_27_Left_139 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_28_Left_140 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_29_Left_141 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_30_Left_142 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_31_Left_143 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_32_Left_144 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_33_Left_145 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_34_Left_146 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_35_Left_147 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_36_Left_148 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_37_Left_149 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_38_Left_150 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_39_Left_151 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_40_Left_152 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_41_Left_153 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_42_Left_154 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_43_Left_155 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_44_Left_156 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_45_Left_157 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_46_Left_158 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_47_Left_159 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_48_Left_160 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_49_Left_161 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_50_Left_162 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_51_Left_163 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_52_Left_164 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_53_Left_165 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_54_Left_166 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_55_Left_167 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_56_Left_168 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_57_Left_169 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_58_Left_170 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_59_Left_171 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_60_Left_172 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_61_Left_173 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_62_Left_174 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_63_Left_175 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_64_Left_176 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_65_Left_177 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_66_Left_178 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_67_Left_179 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_68_Left_180 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_69_Left_181 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_70_Left_182 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_71_Left_183 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_72_Left_184 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_73_Left_185 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_74_Left_186 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_75_Left_187 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_76_Left_188 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_77_Left_189 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_78_Left_190 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_79_Left_191 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_80_Left_192 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_81_Left_193 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_82_Left_194 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_83_Left_195 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_84_Left_196 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_85_Left_197 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_86_Left_198 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_87_Left_199 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_88_Left_200 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_89_Left_201 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_90_Left_202 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_91_Left_203 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_92_Left_204 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_93_Left_205 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_94_Left_206 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_95_Left_207 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_96_Left_208 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_97_Left_209 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_98_Left_210 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_99_Left_211 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_100_Left_212 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_101_Left_213 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_102_Left_214 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_103_Left_215 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_104_Left_216 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_105_Left_217 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_106_Left_218 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_107_Left_219 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_108_Left_220 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_109_Left_221 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_110_Left_222 ();
 sky130_fd_sc_hd__decap_3 PHY_EDGE_ROW_111_Left_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_0_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_1_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_2_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_3_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_4_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_5_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_6_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_7_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_8_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_9_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_10_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_11_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_12_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_13_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_14_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_15_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_16_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_17_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_18_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_19_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_20_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_21_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_22_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_23_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_24_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_25_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_26_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_27_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_28_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_29_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_30_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_31_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_32_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_33_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_34_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_35_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_36_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_37_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_38_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_39_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_40_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_41_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_42_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_43_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_44_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_45_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_46_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_47_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_48_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_49_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_50_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_51_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_52_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_53_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_54_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_55_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_56_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_57_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_58_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_59_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_60_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_61_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_62_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_63_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_64_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_65_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_66_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_67_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_68_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_69_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_70_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_71_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_72_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_73_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_74_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_75_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_76_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_77_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_78_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_79_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_80_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_81_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_82_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_83_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_84_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_85_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_86_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_87_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_88_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_89_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_90_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_91_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_92_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_93_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_94_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_95_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_96_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_97_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_98_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_99_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_100_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_101_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_102_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_103_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_104_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_105_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_106_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_107_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_108_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_109_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_110_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_TAPCELL_ROW_111_1534 ();
endmodule
