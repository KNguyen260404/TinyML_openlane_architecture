module tree_rom_1 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000A43C2154C5000000000110A3;
    rom[1] = 120'h001A43600000C00000000020793;
    rom[2] = 120'h002A4323E9C8700000000030543;
    rom[3] = 120'h003A416FFE2A8000000000402B3;
    rom[4] = 120'h0041406E1000000000000050123;
    rom[5] = 120'h005041D8EC33B00000000060113;
    rom[6] = 120'h006A40CFF7800000000000700C3;
    rom[7] = 120'h007A3FE000000000000000800B3;
    rom[8] = 120'h008041D8EC335000000000900A3;
    rom[9] = 120'h009300000000000000000000001;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00C1406910000000000000D00E3;
    rom[13] = 120'h00D300000000000000000000001;
    rom[14] = 120'h00E1406930000000000000F0103;
    rom[15] = 120'h00F300000000000000000000000;
    rom[16] = 120'h010300000000000000000000001;
    rom[17] = 120'h011300000000000000000000000;
    rom[18] = 120'h0121408A5400000000000130223;
    rom[19] = 120'h0131407F38000000000001401B3;
    rom[20] = 120'h014041D8EC33700000000150183;
    rom[21] = 120'h0151407CC800000000000160173;
    rom[22] = 120'h016300000000000000000000000;
    rom[23] = 120'h017300000000000000000000000;
    rom[24] = 120'h01814077E8000000000001901A3;
    rom[25] = 120'h019300000000000000000000000;
    rom[26] = 120'h01A300000000000000000000000;
    rom[27] = 120'h01BA3FE000000000000001C01F3;
    rom[28] = 120'h01C041D8EC337000000001D01E3;
    rom[29] = 120'h01D300000000000000000000000;
    rom[30] = 120'h01E300000000000000000000000;
    rom[31] = 120'h01F041D8EC33900000000200213;
    rom[32] = 120'h020300000000000000000000001;
    rom[33] = 120'h021300000000000000000000000;
    rom[34] = 120'h022041D8EC339000000002302A3;
    rom[35] = 120'h0231408FDC00000000000240273;
    rom[36] = 120'h024A3FE00000000000000250263;
    rom[37] = 120'h025300000000000000000000000;
    rom[38] = 120'h026300000000000000000000001;
    rom[39] = 120'h027041D8EC33700000000280293;
    rom[40] = 120'h028300000000000000000000001;
    rom[41] = 120'h029300000000000000000000001;
    rom[42] = 120'h02A300000000000000000000000;
    rom[43] = 120'h02B041D8EC33B000000002C04B3;
    rom[44] = 120'h02C041D8EC337000000002D03C3;
    rom[45] = 120'h02D1408A54000000000002E0353;
    rom[46] = 120'h02E041D8EC335000000002F0323;
    rom[47] = 120'h02FA41CA0F72E00000000300313;
    rom[48] = 120'h030300000000000000000000000;
    rom[49] = 120'h031300000000000000000000000;
    rom[50] = 120'h032140680000000000000330343;
    rom[51] = 120'h033300000000000000000000001;
    rom[52] = 120'h034300000000000000000000000;
    rom[53] = 120'h0351409DC200000000000360393;
    rom[54] = 120'h03614093A600000000000370383;
    rom[55] = 120'h037300000000000000000000001;
    rom[56] = 120'h038300000000000000000000001;
    rom[57] = 120'h0391409DCE000000000003A03B3;
    rom[58] = 120'h03A300000000000000000000000;
    rom[59] = 120'h03B300000000000000000000001;
    rom[60] = 120'h03CA41F800000000000003D0443;
    rom[61] = 120'h03D041D8EC339000000003E0413;
    rom[62] = 120'h03E1408A5C000000000003F0403;
    rom[63] = 120'h03F300000000000000000000000;
    rom[64] = 120'h040300000000000000000000001;
    rom[65] = 120'h041A41EFF150000000000420433;
    rom[66] = 120'h042300000000000000000000000;
    rom[67] = 120'h043300000000000000000000001;
    rom[68] = 120'h044140783800000000000450483;
    rom[69] = 120'h045A42D00000200000000460473;
    rom[70] = 120'h046300000000000000000000001;
    rom[71] = 120'h047300000000000000000000000;
    rom[72] = 120'h048A4313EC584000000004904A3;
    rom[73] = 120'h049300000000000000000000000;
    rom[74] = 120'h04A300000000000000000000000;
    rom[75] = 120'h04BA421C00000000000004C04D3;
    rom[76] = 120'h04C300000000000000000000000;
    rom[77] = 120'h04D1408B88000000000004E04F3;
    rom[78] = 120'h04E300000000000000000000000;
    rom[79] = 120'h04F1408F8800000000000500533;
    rom[80] = 120'h050A42755000000000000510523;
    rom[81] = 120'h051300000000000000000000001;
    rom[82] = 120'h052300000000000000000000000;
    rom[83] = 120'h053300000000000000000000000;
    rom[84] = 120'h054A432400181000000005505E3;
    rom[85] = 120'h055041D8EC339000000005605D3;
    rom[86] = 120'h056041D8EC33500000000570583;
    rom[87] = 120'h057300000000000000000000001;
    rom[88] = 120'h058041D8EC337000000005905A3;
    rom[89] = 120'h059300000000000000000000001;
    rom[90] = 120'h05A1408990000000000005B05C3;
    rom[91] = 120'h05B300000000000000000000001;
    rom[92] = 120'h05C300000000000000000000001;
    rom[93] = 120'h05D300000000000000000000000;
    rom[94] = 120'h05E041D8EC339000000005F0783;
    rom[95] = 120'h05F14068D0000000000006006B3;
    rom[96] = 120'h060A434DD445A00000000610663;
    rom[97] = 120'h061A432684B3500000000620633;
    rom[98] = 120'h062300000000000000000000000;
    rom[99] = 120'h063041D8EC33700000000640653;
    rom[100] = 120'h064300000000000000000000001;
    rom[101] = 120'h065300000000000000000000000;
    rom[102] = 120'h066140681000000000000670683;
    rom[103] = 120'h067300000000000000000000001;
    rom[104] = 120'h068A434F1C26C000000006906A3;
    rom[105] = 120'h069300000000000000000000000;
    rom[106] = 120'h06A300000000000000000000000;
    rom[107] = 120'h06B1407E88000000000006C0713;
    rom[108] = 120'h06C041D8EC335000000006D0703;
    rom[109] = 120'h06D1406940000000000006E06F3;
    rom[110] = 120'h06E300000000000000000000000;
    rom[111] = 120'h06F300000000000000000000001;
    rom[112] = 120'h070300000000000000000000001;
    rom[113] = 120'h071041D8EC33700000000720753;
    rom[114] = 120'h0721407E9800000000000730743;
    rom[115] = 120'h073300000000000000000000000;
    rom[116] = 120'h074300000000000000000000001;
    rom[117] = 120'h075A43565894900000000760773;
    rom[118] = 120'h076300000000000000000000000;
    rom[119] = 120'h077300000000000000000000001;
    rom[120] = 120'h078300000000000000000000000;
    rom[121] = 120'h0791407E98000000000007A0CB3;
    rom[122] = 120'h07AA43700192F000000007B09C3;
    rom[123] = 120'h07B041D8EC337000000007C0933;
    rom[124] = 120'h07CA4360815FC000000007D08A3;
    rom[125] = 120'h07D041D8EC335000000007E0853;
    rom[126] = 120'h07E1406B70000000000007F0823;
    rom[127] = 120'h07F14065B000000000000800813;
    rom[128] = 120'h080300000000000000000000001;
    rom[129] = 120'h081300000000000000000000000;
    rom[130] = 120'h0821407BD800000000000830843;
    rom[131] = 120'h083300000000000000000000001;
    rom[132] = 120'h084300000000000000000000000;
    rom[133] = 120'h085A436014CFE00000000860873;
    rom[134] = 120'h086300000000000000000000000;
    rom[135] = 120'h0871406FB000000000000880893;
    rom[136] = 120'h088300000000000000000000000;
    rom[137] = 120'h089300000000000000000000001;
    rom[138] = 120'h08AA436081603000000008B08C3;
    rom[139] = 120'h08B300000000000000000000001;
    rom[140] = 120'h08C041D8EC335000000008D0903;
    rom[141] = 120'h08DA436089922000000008E08F3;
    rom[142] = 120'h08E300000000000000000000000;
    rom[143] = 120'h08F300000000000000000000001;
    rom[144] = 120'h090A43700052800000000910923;
    rom[145] = 120'h091300000000000000000000000;
    rom[146] = 120'h092300000000000000000000001;
    rom[147] = 120'h093A43600600200000000940953;
    rom[148] = 120'h094300000000000000000000000;
    rom[149] = 120'h095A43600A52800000000960973;
    rom[150] = 120'h096300000000000000000000001;
    rom[151] = 120'h097140680000000000000980993;
    rom[152] = 120'h098300000000000000000000001;
    rom[153] = 120'h099A436FEAACA000000009A09B3;
    rom[154] = 120'h09A300000000000000000000000;
    rom[155] = 120'h09B300000000000000000000000;
    rom[156] = 120'h09CA43B400D0F000000009D0B43;
    rom[157] = 120'h09D041D8EC337000000009E0A73;
    rom[158] = 120'h09E1406810000000000009F0A03;
    rom[159] = 120'h09F300000000000000000000001;
    rom[160] = 120'h0A0041D8EC33500000000A10A43;
    rom[161] = 120'h0A114068F000000000000A20A33;
    rom[162] = 120'h0A2300000000000000000000000;
    rom[163] = 120'h0A3300000000000000000000000;
    rom[164] = 120'h0A414077C000000000000A50A63;
    rom[165] = 120'h0A5300000000000000000000000;
    rom[166] = 120'h0A6300000000000000000000000;
    rom[167] = 120'h0A7A43A04899300000000A80AF3;
    rom[168] = 120'h0A8A4399D659400000000A90AC3;
    rom[169] = 120'h0A9041D8EC33900000000AA0AB3;
    rom[170] = 120'h0AA300000000000000000000000;
    rom[171] = 120'h0AB300000000000000000000000;
    rom[172] = 120'h0ACA439A8439E00000000AD0AE3;
    rom[173] = 120'h0AD300000000000000000000000;
    rom[174] = 120'h0AE300000000000000000000000;
    rom[175] = 120'h0AF041D8EC33900000000B00B33;
    rom[176] = 120'h0B0140673000000000000B10B23;
    rom[177] = 120'h0B1300000000000000000000001;
    rom[178] = 120'h0B2300000000000000000000000;
    rom[179] = 120'h0B3300000000000000000000000;
    rom[180] = 120'h0B4041D8EC33700000000B50C43;
    rom[181] = 120'h0B5041D8EC33500000000B60BD3;
    rom[182] = 120'h0B6A43BFFF45300000000B70BA3;
    rom[183] = 120'h0B7140798800000000000B80B93;
    rom[184] = 120'h0B8300000000000000000000001;
    rom[185] = 120'h0B9300000000000000000000001;
    rom[186] = 120'h0BA14068C000000000000BB0BC3;
    rom[187] = 120'h0BB300000000000000000000000;
    rom[188] = 120'h0BC300000000000000000000001;
    rom[189] = 120'h0BD14068B000000000000BE0C13;
    rom[190] = 120'h0BEA43BFF8BCB00000000BF0C03;
    rom[191] = 120'h0BF300000000000000000000001;
    rom[192] = 120'h0C0300000000000000000000000;
    rom[193] = 120'h0C1A43B84BD4800000000C20C33;
    rom[194] = 120'h0C2300000000000000000000001;
    rom[195] = 120'h0C3300000000000000000000001;
    rom[196] = 120'h0C4041D8EC33900000000C50CA3;
    rom[197] = 120'h0C514066E000000000000C60C73;
    rom[198] = 120'h0C6300000000000000000000001;
    rom[199] = 120'h0C71406B2000000000000C80C93;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C9300000000000000000000001;
    rom[202] = 120'h0CA300000000000000000000000;
    rom[203] = 120'h0CBA43A00BD3A00000000CC0E73;
    rom[204] = 120'h0CC14093C800000000000CD0E63;
    rom[205] = 120'h0CD1407F6800000000000CE0D93;
    rom[206] = 120'h0CE041D8EC33500000000CF0D43;
    rom[207] = 120'h0CFA436D9295E00000000D00D13;
    rom[208] = 120'h0D0300000000000000000000001;
    rom[209] = 120'h0D1A439036C4380000000D20D33;
    rom[210] = 120'h0D2300000000000000000000000;
    rom[211] = 120'h0D3300000000000000000000001;
    rom[212] = 120'h0D41407F4800000000000D50D63;
    rom[213] = 120'h0D5300000000000000000000001;
    rom[214] = 120'h0D6A436CDD0CC00000000D70D83;
    rom[215] = 120'h0D7300000000000000000000001;
    rom[216] = 120'h0D8300000000000000000000000;
    rom[217] = 120'h0D9041D8EC33700000000DA0E13;
    rom[218] = 120'h0DAA439D93B0A00000000DB0DE3;
    rom[219] = 120'h0DB041D8EC33500000000DC0DD3;
    rom[220] = 120'h0DC300000000000000000000001;
    rom[221] = 120'h0DD300000000000000000000001;
    rom[222] = 120'h0DE1408D9800000000000DF0E03;
    rom[223] = 120'h0DF300000000000000000000001;
    rom[224] = 120'h0E0300000000000000000000000;
    rom[225] = 120'h0E1041D8EC33900000000E20E53;
    rom[226] = 120'h0E2A436A0D7A200000000E30E43;
    rom[227] = 120'h0E3300000000000000000000001;
    rom[228] = 120'h0E4300000000000000000000000;
    rom[229] = 120'h0E5300000000000000000000000;
    rom[230] = 120'h0E6300000000000000000000001;
    rom[231] = 120'h0E7A43C201FAA00000000E81033;
    rom[232] = 120'h0E81408F4000000000000E90F63;
    rom[233] = 120'h0E9041D8EC33900000000EA0F13;
    rom[234] = 120'h0EA041D8EC33500000000EB0EE3;
    rom[235] = 120'h0EBA43AE7564100000000EC0ED3;
    rom[236] = 120'h0EC300000000000000000000000;
    rom[237] = 120'h0ED300000000000000000000001;
    rom[238] = 120'h0EE1407F6000000000000EF0F03;
    rom[239] = 120'h0EF300000000000000000000001;
    rom[240] = 120'h0F0300000000000000000000001;
    rom[241] = 120'h0F1041D8EC33B00000000F20F53;
    rom[242] = 120'h0F2A43AB1B00000000000F30F43;
    rom[243] = 120'h0F3300000000000000000000001;
    rom[244] = 120'h0F4300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule

