module tree_rom_15 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000140681000000000000010023;
    rom[1] = 120'h001300000000000000000000001;
    rom[2] = 120'h002A43D3FFE4D00000000030A43;
    rom[3] = 120'h003041D8EC339000000000407F3;
    rom[4] = 120'h004A4360009C400000000050423;
    rom[5] = 120'h005041D8EC33500000000060233;
    rom[6] = 120'h006A4170180BC00000000070143;
    rom[7] = 120'h007A41391EFA0000000000800F3;
    rom[8] = 120'h0081406890000000000000900C3;
    rom[9] = 120'h0091406830000000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000001;
    rom[12] = 120'h00CA3FE000000000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000001;
    rom[15] = 120'h00F1408A5800000000000100133;
    rom[16] = 120'h010A4162B27C900000000110123;
    rom[17] = 120'h011300000000000000000000001;
    rom[18] = 120'h012300000000000000000000001;
    rom[19] = 120'h013300000000000000000000001;
    rom[20] = 120'h014A4322F78B7000000001501C3;
    rom[21] = 120'h0151408A5400000000000160193;
    rom[22] = 120'h016A41D2AD96500000000170183;
    rom[23] = 120'h017300000000000000000000000;
    rom[24] = 120'h018300000000000000000000000;
    rom[25] = 120'h01914093A6000000000001A01B3;
    rom[26] = 120'h01A300000000000000000000001;
    rom[27] = 120'h01B300000000000000000000001;
    rom[28] = 120'h01CA432400181000000001D0203;
    rom[29] = 120'h01D1407FE8000000000001E01F3;
    rom[30] = 120'h01E300000000000000000000001;
    rom[31] = 120'h01F300000000000000000000001;
    rom[32] = 120'h020A435269E8B00000000210223;
    rom[33] = 120'h021300000000000000000000001;
    rom[34] = 120'h022300000000000000000000001;
    rom[35] = 120'h0231408A5400000000000240333;
    rom[36] = 120'h024A4322C8C43000000002502C3;
    rom[37] = 120'h025041D8EC33700000000260293;
    rom[38] = 120'h026A40040000000000000270283;
    rom[39] = 120'h027300000000000000000000000;
    rom[40] = 120'h028300000000000000000000000;
    rom[41] = 120'h0291406E10000000000002A02B3;
    rom[42] = 120'h02A300000000000000000000001;
    rom[43] = 120'h02B300000000000000000000000;
    rom[44] = 120'h02CA432400181000000002D0303;
    rom[45] = 120'h02DA4323CDB21000000002E02F3;
    rom[46] = 120'h02E300000000000000000000001;
    rom[47] = 120'h02F300000000000000000000001;
    rom[48] = 120'h03014068D000000000000310323;
    rom[49] = 120'h031300000000000000000000000;
    rom[50] = 120'h032300000000000000000000001;
    rom[51] = 120'h0331408FC4000000000003403B3;
    rom[52] = 120'h034041D8EC33700000000350383;
    rom[53] = 120'h035A3FE00000000000000360373;
    rom[54] = 120'h036300000000000000000000000;
    rom[55] = 120'h037300000000000000000000001;
    rom[56] = 120'h038A4278A3FCA000000003903A3;
    rom[57] = 120'h039300000000000000000000001;
    rom[58] = 120'h03A300000000000000000000001;
    rom[59] = 120'h03BA3FE000000000000003C03F3;
    rom[60] = 120'h03C14093B4000000000003D03E3;
    rom[61] = 120'h03D300000000000000000000000;
    rom[62] = 120'h03E300000000000000000000000;
    rom[63] = 120'h03F041D8EC33700000000400413;
    rom[64] = 120'h040300000000000000000000001;
    rom[65] = 120'h041300000000000000000000001;
    rom[66] = 120'h042A43A0B45D500000000430623;
    rom[67] = 120'h0431407F6000000000000440533;
    rom[68] = 120'h044A437002BB1000000004504C3;
    rom[69] = 120'h0451406F3000000000000460493;
    rom[70] = 120'h046A43600720800000000470483;
    rom[71] = 120'h047300000000000000000000000;
    rom[72] = 120'h048300000000000000000000000;
    rom[73] = 120'h049A436BA0E78000000004A04B3;
    rom[74] = 120'h04A300000000000000000000001;
    rom[75] = 120'h04B300000000000000000000001;
    rom[76] = 120'h04C1407900000000000004D0503;
    rom[77] = 120'h04D1406F60000000000004E04F3;
    rom[78] = 120'h04E300000000000000000000000;
    rom[79] = 120'h04F300000000000000000000000;
    rom[80] = 120'h050A4397FE2F400000000510523;
    rom[81] = 120'h051300000000000000000000000;
    rom[82] = 120'h052300000000000000000000000;
    rom[83] = 120'h053A439D93B0A000000005405B3;
    rom[84] = 120'h054A436FEB0F400000000550583;
    rom[85] = 120'h055140930A00000000000560573;
    rom[86] = 120'h056300000000000000000000001;
    rom[87] = 120'h057300000000000000000000001;
    rom[88] = 120'h05814093D0000000000005905A3;
    rom[89] = 120'h059300000000000000000000001;
    rom[90] = 120'h05A300000000000000000000001;
    rom[91] = 120'h05B041D8EC337000000005C05F3;
    rom[92] = 120'h05C041D8EC335000000005D05E3;
    rom[93] = 120'h05D300000000000000000000000;
    rom[94] = 120'h05E300000000000000000000000;
    rom[95] = 120'h05F1408BF400000000000600613;
    rom[96] = 120'h060300000000000000000000001;
    rom[97] = 120'h061300000000000000000000000;
    rom[98] = 120'h0621407E9800000000000630703;
    rom[99] = 120'h063A43ADD5A7200000000640693;
    rom[100] = 120'h064140790800000000000650663;
    rom[101] = 120'h065300000000000000000000001;
    rom[102] = 120'h066A43A1E558100000000670683;
    rom[103] = 120'h067300000000000000000000000;
    rom[104] = 120'h068300000000000000000000001;
    rom[105] = 120'h069041D8EC337000000006A06D3;
    rom[106] = 120'h06AA43D17E79E000000006B06C3;
    rom[107] = 120'h06B300000000000000000000000;
    rom[108] = 120'h06C300000000000000000000000;
    rom[109] = 120'h06DA43D17BE98000000006E06F3;
    rom[110] = 120'h06E300000000000000000000000;
    rom[111] = 120'h06F300000000000000000000000;
    rom[112] = 120'h070A43AB734B400000000710783;
    rom[113] = 120'h071A43A96B89C00000000720753;
    rom[114] = 120'h072041D8EC33700000000730743;
    rom[115] = 120'h073300000000000000000000001;
    rom[116] = 120'h074300000000000000000000001;
    rom[117] = 120'h075041D8EC33700000000760773;
    rom[118] = 120'h076300000000000000000000001;
    rom[119] = 120'h077300000000000000000000001;
    rom[120] = 120'h078041D8EC335000000007907C3;
    rom[121] = 120'h0791407F58000000000007A07B3;
    rom[122] = 120'h07A300000000000000000000000;
    rom[123] = 120'h07B300000000000000000000001;
    rom[124] = 120'h07CA43AE1E002000000007D07E3;
    rom[125] = 120'h07D300000000000000000000000;
    rom[126] = 120'h07E300000000000000000000001;
    rom[127] = 120'h07F1408EE800000000000800973;
    rom[128] = 120'h080041D8EC33B00000000810963;
    rom[129] = 120'h0811406BA000000000000820893;
    rom[130] = 120'h082A419C0082100000000830883;
    rom[131] = 120'h083A40C00800000000000840853;
    rom[132] = 120'h084300000000000000000000001;
    rom[133] = 120'h085A418C0104200000000860873;
    rom[134] = 120'h086300000000000000000000000;
    rom[135] = 120'h087300000000000000000000001;
    rom[136] = 120'h088300000000000000000000000;
    rom[137] = 120'h089A42D000002000000008A0913;
    rom[138] = 120'h08A14075F8000000000008B08E3;
    rom[139] = 120'h08BA42C0002ECF80000008C08D3;
    rom[140] = 120'h08C300000000000000000000000;
    rom[141] = 120'h08D300000000000000000000001;
    rom[142] = 120'h08EA420D9010E000000008F0903;
    rom[143] = 120'h08F300000000000000000000000;
    rom[144] = 120'h090300000000000000000000000;
    rom[145] = 120'h0911407EF000000000000920933;
    rom[146] = 120'h092300000000000000000000000;
    rom[147] = 120'h093A43A47300000000000940953;
    rom[148] = 120'h094300000000000000000000000;
    rom[149] = 120'h095300000000000000000000000;
    rom[150] = 120'h096300000000000000000000000;
    rom[151] = 120'h097A425D680B8000000009809D3;
    rom[152] = 120'h0981408F90000000000009909C3;
    rom[153] = 120'h099A41E000000000000009A09B3;
    rom[154] = 120'h09A300000000000000000000000;
    rom[155] = 120'h09B300000000000000000000001;
    rom[156] = 120'h09C300000000000000000000000;
    rom[157] = 120'h09D041D8EC33D000000009E0A33;
    rom[158] = 120'h09E1408F68000000000009F0A23;
    rom[159] = 120'h09FA43BBF184C00000000A00A13;
    rom[160] = 120'h0A0300000000000000000000000;
    rom[161] = 120'h0A1300000000000000000000001;
    rom[162] = 120'h0A2300000000000000000000000;
    rom[163] = 120'h0A3300000000000000000000000;
    rom[164] = 120'h0A4041D8EC33900000000A50E63;
    rom[165] = 120'h0A51407F1800000000000A60D73;
    rom[166] = 120'h0A6041D8EC33500000000A70C23;
    rom[167] = 120'h0A7140798800000000000A80B33;
    rom[168] = 120'h0A81406F3000000000000A90AE3;
    rom[169] = 120'h0A9A43DF7718D00000000AA0AD3;
    rom[170] = 120'h0AA1406F1000000000000AB0AC3;
    rom[171] = 120'h0AB300000000000000000000001;
    rom[172] = 120'h0AC300000000000000000000000;
    rom[173] = 120'h0AD300000000000000000000001;
    rom[174] = 120'h0AEA43D5BBBD700000000AF0B03;
    rom[175] = 120'h0AF300000000000000000000001;
    rom[176] = 120'h0B0A43D5C3A9F00000000B10B23;
    rom[177] = 120'h0B1300000000000000000000000;
    rom[178] = 120'h0B2300000000000000000000001;
    rom[179] = 120'h0B314079D800000000000B40BB3;
    rom[180] = 120'h0B4140799800000000000B50B83;
    rom[181] = 120'h0B5A43E05597880000000B60B73;
    rom[182] = 120'h0B6300000000000000000000001;
    rom[183] = 120'h0B7300000000000000000000000;
    rom[184] = 120'h0B8A43EC4978200000000B90BA3;
    rom[185] = 120'h0B9300000000000000000000000;
    rom[186] = 120'h0BA300000000000000000000001;
    rom[187] = 120'h0BBA43E5C750700000000BC0BF3;
    rom[188] = 120'h0BC1407F0800000000000BD0BE3;
    rom[189] = 120'h0BD300000000000000000000001;
    rom[190] = 120'h0BE300000000000000000000000;
    rom[191] = 120'h0BFA43E76255000000000C00C13;
    rom[192] = 120'h0C0300000000000000000000001;
    rom[193] = 120'h0C1300000000000000000000001;
    rom[194] = 120'h0C2041D8EC33700000000C30D03;
    rom[195] = 120'h0C3A43DFFC0A000000000C40C93;
    rom[196] = 120'h0C4A43D5F6CA500000000C50C83;
    rom[197] = 120'h0C5140796800000000000C60C73;
    rom[198] = 120'h0C6300000000000000000000001;
    rom[199] = 120'h0C7300000000000000000000001;
    rom[200] = 120'h0C8300000000000000000000001;
    rom[201] = 120'h0C9A43EA02F4500000000CA0CD3;
    rom[202] = 120'h0CAA43E9FCB0200000000CB0CC3;
    rom[203] = 120'h0CB300000000000000000000000;
    rom[204] = 120'h0CC300000000000000000000000;
    rom[205] = 120'h0CDA43EAFD57800000000CE0CF3;
    rom[206] = 120'h0CE300000000000000000000001;
    rom[207] = 120'h0CF300000000000000000000001;
    rom[208] = 120'h0D0140798000000000000D10D23;
    rom[209] = 120'h0D1300000000000000000000001;
    rom[210] = 120'h0D2A43EA163C600000000D30D63;
    rom[211] = 120'h0D314079E800000000000D40D53;
    rom[212] = 120'h0D4300000000000000000000000;
    rom[213] = 120'h0D5300000000000000000000000;
    rom[214] = 120'h0D6300000000000000000000001;
    rom[215] = 120'h0D7A43E00094B00000000D80E53;
    rom[216] = 120'h0D8041D8EC33700000000D90E23;
    rom[217] = 120'h0D9041D8EC33500000000DA0DD3;
    rom[218] = 120'h0DAA43DFFF61A00000000DB0DC3;
    rom[219] = 120'h0DB300000000000000000000001;
    rom[220] = 120'h0DC300000000000000000000000;
    rom[221] = 120'h0DD1408F7000000000000DE0E13;
    rom[222] = 120'h0DE1408F6000000000000DF0E03;
    rom[223] = 120'h0DF300000000000000000000001;
    rom[224] = 120'h0E0300000000000000000000000;
    rom[225] = 120'h0E1300000000000000000000001;
    rom[226] = 120'h0E2A43DFFD1AF00000000E30E43;
    rom[227] = 120'h0E3300000000000000000000001;
    rom[228] = 120'h0E4300000000000000000000000;
    rom[229] = 120'h0E5300000000000000000000001;
    rom[230] = 120'h0E6300000000000000000000000;
    // Initialize remaining locations with zeros
    for (integer i = 231; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 

