module tree_rom_6 #(
    parameter NODE_WIDTH = 120,
    parameter ADDR_WIDTH = 10,
    parameter ROM_DEPTH = 512
)(
    input wire clk,
    input wire [ADDR_WIDTH-1:0] addr,
    output reg [NODE_WIDTH-1:0] node_data
);

reg [NODE_WIDTH-1:0] rom [0:ROM_DEPTH-1];

// Define a 9-bit address for properly indexing into the ROM
wire [8:0] rom_addr = addr[8:0];

initial begin
    rom[0] = 120'h000140681000000000000010023;
    rom[1] = 120'h001300000000000000000000001;
    rom[2] = 120'h002A43D3FFCBB00000000030A63;
    rom[3] = 120'h003A43600000C000000000405D3;
    rom[4] = 120'h0041408A54000000000000503C3;
    rom[5] = 120'h005A4323ED19000000000060233;
    rom[6] = 120'h0061406E1000000000000070143;
    rom[7] = 120'h0071406890000000000000800F3;
    rom[8] = 120'h008A4203FB67E000000000900C3;
    rom[9] = 120'h009041D8EC335000000000A00B3;
    rom[10] = 120'h00A300000000000000000000001;
    rom[11] = 120'h00B300000000000000000000000;
    rom[12] = 120'h00C041D8EC335000000000D00E3;
    rom[13] = 120'h00D300000000000000000000000;
    rom[14] = 120'h00E300000000000000000000000;
    rom[15] = 120'h00F041D8EC33B00000000100133;
    rom[16] = 120'h010041D8EC33700000000110123;
    rom[17] = 120'h011300000000000000000000001;
    rom[18] = 120'h012300000000000000000000001;
    rom[19] = 120'h013300000000000000000000000;
    rom[20] = 120'h0141407F38000000000001501C3;
    rom[21] = 120'h015041D8EC33700000000160193;
    rom[22] = 120'h016A40040000000000000170183;
    rom[23] = 120'h017300000000000000000000000;
    rom[24] = 120'h018300000000000000000000000;
    rom[25] = 120'h019041D8EC33B000000001A01B3;
    rom[26] = 120'h01A300000000000000000000000;
    rom[27] = 120'h01B300000000000000000000000;
    rom[28] = 120'h01C041D8EC337000000001D0203;
    rom[29] = 120'h01D041D8EC335000000001E01F3;
    rom[30] = 120'h01E300000000000000000000001;
    rom[31] = 120'h01F300000000000000000000000;
    rom[32] = 120'h020140861400000000000210223;
    rom[33] = 120'h021300000000000000000000001;
    rom[34] = 120'h022300000000000000000000000;
    rom[35] = 120'h02314068D000000000000240313;
    rom[36] = 120'h024A435E504DF000000002502C3;
    rom[37] = 120'h025A433DD9C7900000000260293;
    rom[38] = 120'h026041D8EC33700000000270283;
    rom[39] = 120'h027300000000000000000000000;
    rom[40] = 120'h028300000000000000000000000;
    rom[41] = 120'h029041D8EC337000000002A02B3;
    rom[42] = 120'h02A300000000000000000000000;
    rom[43] = 120'h02B300000000000000000000000;
    rom[44] = 120'h02C1406850000000000002D02E3;
    rom[45] = 120'h02D300000000000000000000000;
    rom[46] = 120'h02E1406890000000000002F0303;
    rom[47] = 120'h02F300000000000000000000001;
    rom[48] = 120'h030300000000000000000000000;
    rom[49] = 120'h031A43240018100000000320373;
    rom[50] = 120'h032041D8EC33900000000330363;
    rom[51] = 120'h033041D8EC33700000000340353;
    rom[52] = 120'h034300000000000000000000001;
    rom[53] = 120'h035300000000000000000000001;
    rom[54] = 120'h036300000000000000000000000;
    rom[55] = 120'h037041D8EC339000000003803B3;
    rom[56] = 120'h0381407E78000000000003903A3;
    rom[57] = 120'h039300000000000000000000001;
    rom[58] = 120'h03A300000000000000000000001;
    rom[59] = 120'h03B300000000000000000000000;
    rom[60] = 120'h03C1409DC2000000000003D0523;
    rom[61] = 120'h03DA3FE000000000000003E0453;
    rom[62] = 120'h03E041D8EC337000000003F0443;
    rom[63] = 120'h03F140943600000000000400433;
    rom[64] = 120'h0401408ED400000000000410423;
    rom[65] = 120'h041300000000000000000000001;
    rom[66] = 120'h042300000000000000000000000;
    rom[67] = 120'h043300000000000000000000001;
    rom[68] = 120'h044300000000000000000000000;
    rom[69] = 120'h045A426C2450F000000004604D3;
    rom[70] = 120'h046A40838C000000000004704A3;
    rom[71] = 120'h0471408FE000000000000480493;
    rom[72] = 120'h048300000000000000000000000;
    rom[73] = 120'h049300000000000000000000001;
    rom[74] = 120'h04AA41D681A5D000000004B04C3;
    rom[75] = 120'h04B300000000000000000000001;
    rom[76] = 120'h04C300000000000000000000001;
    rom[77] = 120'h04DA426C28161000000004E04F3;
    rom[78] = 120'h04E300000000000000000000000;
    rom[79] = 120'h04F1408FCC00000000000500513;
    rom[80] = 120'h050300000000000000000000000;
    rom[81] = 120'h051300000000000000000000001;
    rom[82] = 120'h052A3FE00000000000000530543;
    rom[83] = 120'h053300000000000000000000000;
    rom[84] = 120'h054041D8EC339000000005505C3;
    rom[85] = 120'h055A42C3C1205D00000000560593;
    rom[86] = 120'h056A42B0C5C2100000000570583;
    rom[87] = 120'h057300000000000000000000001;
    rom[88] = 120'h058300000000000000000000001;
    rom[89] = 120'h0591409DCE000000000005A05B3;
    rom[90] = 120'h05A300000000000000000000000;
    rom[91] = 120'h05B300000000000000000000001;
    rom[92] = 120'h05C300000000000000000000000;
    rom[93] = 120'h05D041D8EC339000000005E09B3;
    rom[94] = 120'h05E041D8EC337000000005F07E3;
    rom[95] = 120'h05F1407E98000000000006006F3;
    rom[96] = 120'h06014068B000000000000610683;
    rom[97] = 120'h061140683000000000000620653;
    rom[98] = 120'h062A43C9D283300000000630643;
    rom[99] = 120'h063300000000000000000000000;
    rom[100] = 120'h064300000000000000000000000;
    rom[101] = 120'h065041D8EC33500000000660673;
    rom[102] = 120'h066300000000000000000000000;
    rom[103] = 120'h067300000000000000000000000;
    rom[104] = 120'h0681407908000000000006906C3;
    rom[105] = 120'h069A431207ED44000000006A06B3;
    rom[106] = 120'h06A300000000000000000000000;
    rom[107] = 120'h06B300000000000000000000001;
    rom[108] = 120'h06C041D8EC335000000006D06E3;
    rom[109] = 120'h06D300000000000000000000000;
    rom[110] = 120'h06E300000000000000000000000;
    rom[111] = 120'h06FA43A009CD300000000700773;
    rom[112] = 120'h070041D8EC33500000000710743;
    rom[113] = 120'h071A436FEB0F400000000720733;
    rom[114] = 120'h072300000000000000000000001;
    rom[115] = 120'h073300000000000000000000000;
    rom[116] = 120'h074A4374B000000000000750763;
    rom[117] = 120'h075300000000000000000000001;
    rom[118] = 120'h076300000000000000000000000;
    rom[119] = 120'h077A43B2D27B1000000007807B3;
    rom[120] = 120'h0781409308000000000007907A3;
    rom[121] = 120'h079300000000000000000000001;
    rom[122] = 120'h07A300000000000000000000001;
    rom[123] = 120'h07BA43D007FE7000000007C07D3;
    rom[124] = 120'h07C300000000000000000000001;
    rom[125] = 120'h07D300000000000000000000001;
    rom[126] = 120'h07E1407E98000000000007F08E3;
    rom[127] = 120'h07F140790800000000000800873;
    rom[128] = 120'h080A43C2A1E8A00000000810843;
    rom[129] = 120'h08114077E800000000000820833;
    rom[130] = 120'h082300000000000000000000000;
    rom[131] = 120'h083300000000000000000000001;
    rom[132] = 120'h08414072A800000000000850863;
    rom[133] = 120'h085300000000000000000000000;
    rom[134] = 120'h086300000000000000000000001;
    rom[135] = 120'h0871407E48000000000008808B3;
    rom[136] = 120'h0881407C38000000000008908A3;
    rom[137] = 120'h089300000000000000000000000;
    rom[138] = 120'h08A300000000000000000000001;
    rom[139] = 120'h08B1407E60000000000008C08D3;
    rom[140] = 120'h08C300000000000000000000000;
    rom[141] = 120'h08D300000000000000000000000;
    rom[142] = 120'h08EA43A1AB551000000008F0943;
    rom[143] = 120'h08F14093F600000000000900933;
    rom[144] = 120'h0901408F9800000000000910923;
    rom[145] = 120'h091300000000000000000000000;
    rom[146] = 120'h092300000000000000000000000;
    rom[147] = 120'h093300000000000000000000001;
    rom[148] = 120'h094140930000000000000950983;
    rom[149] = 120'h095A43D0F17AA000000001200973;
    rom[150] = 120'h0120300000000000000000000001;
    rom[151] = 120'h097300000000000000000000000;
    rom[152] = 120'h098A43D008641000000009909A3;
    rom[153] = 120'h099300000000000000000000001;
    rom[154] = 120'h09A300000000000000000000000;
    rom[155] = 120'h09BA43AA19180000000009C09D3;
    rom[156] = 120'h09C300000000000000000000000;
    rom[157] = 120'h09D1407EF0000000000009E09F3;
    rom[158] = 120'h09E300000000000000000000000;
    rom[159] = 120'h09FA43AA1B17F00000000A00A13;
    rom[160] = 120'h0A0300000000000000000000001;
    rom[161] = 120'h0A1140877800000000000A20A33;
    rom[162] = 120'h0A2300000000000000000000000;
    rom[163] = 120'h0A3140915400000000000A40A53;
    rom[164] = 120'h0A4300000000000000000000000;
    rom[165] = 120'h0A5300000000000000000000000;
    rom[166] = 120'h0A61407F1800000000000A70EA3;
    rom[167] = 120'h0A7041D8EC33700000000A80D53;
    rom[168] = 120'h0A8041D8EC33500000000A90C23;
    rom[169] = 120'h0A9140798800000000000AA0B53;
    rom[170] = 120'h0AAA43DEC150A00000000AB0B03;
    rom[171] = 120'h0ABA43D5BBBD700000000AC0AD3;
    rom[172] = 120'h0AC300000000000000000000001;
    rom[173] = 120'h0AD140729800000000000AE0AF3;
    rom[174] = 120'h0AE300000000000000000000001;
    rom[175] = 120'h0AF300000000000000000000001;
    rom[176] = 120'h0B01406F3000000000000B10B43;
    rom[177] = 120'h0B11406F1000000000000B20B33;
    rom[178] = 120'h0B2300000000000000000000001;
    rom[179] = 120'h0B3300000000000000000000000;
    rom[180] = 120'h0B4300000000000000000000001;
    rom[181] = 120'h0B5A43EA3BB6300000000B60BD3;
    rom[182] = 120'h0B6A43DFF74E900000000B70BA3;
    rom[183] = 120'h0B7A43D4734A100000000B80B93;
    rom[184] = 120'h0B8300000000000000000000000;
    rom[185] = 120'h0B9300000000000000000000001;
    rom[186] = 120'h0BA14079D800000000000BB0BC3;
    rom[187] = 120'h0BB300000000000000000000000;
    rom[188] = 120'h0BC300000000000000000000001;
    rom[189] = 120'h0BDA43EB0072B00000000BE0C13;
    rom[190] = 120'h0BE14079A800000000000BF0C03;
    rom[191] = 120'h0BF300000000000000000000000;
    rom[192] = 120'h0C0300000000000000000000001;
    rom[193] = 120'h0C1300000000000000000000001;
    rom[194] = 120'h0C2A43DFFC0A000000000C30CA3;
    rom[195] = 120'h0C3A43D5F772400000000C40C93;
    rom[196] = 120'h0C4A43D5C44FF00000000C50C63;
    rom[197] = 120'h0C5300000000000000000000001;
    rom[198] = 120'h0C614077F000000000000C70C83;
    rom[199] = 120'h0C7300000000000000000000001;
    rom[200] = 120'h0C8300000000000000000000000;
    rom[201] = 120'h0C9300000000000000000000001;
    rom[202] = 120'h0CAA43EA007B200000000CB0D03;
    rom[203] = 120'h0CBA43E9FCB0200000000CC0CF3;
    rom[204] = 120'h0CCA43E20011B00000000CD0CE3;
    rom[205] = 120'h0CD300000000000000000000000;
    rom[206] = 120'h0CE300000000000000000000001;
    rom[207] = 120'h0CF300000000000000000000000;
    rom[208] = 120'h0D0140798800000000000D10D23;
    rom[209] = 120'h0D1300000000000000000000001;
    rom[210] = 120'h0D2140799800000000000D30D43;
    rom[211] = 120'h0D3300000000000000000000000;
    rom[212] = 120'h0D4300000000000000000000001;
    rom[213] = 120'h0D5140798000000000000D60D93;
    rom[214] = 120'h0D6041D8EC33900000000D70D83;
    rom[215] = 120'h0D7300000000000000000000001;
    rom[216] = 120'h0D8300000000000000000000000;
    rom[217] = 120'h0D9A43EA163C600000000DA0E33;
    rom[218] = 120'h0DA041D8EC33900000000DB0E23;
    rom[219] = 120'h0DBA43DFDE11200000000DC0DF3;
    rom[220] = 120'h0DCA43D60E23500000000DD0DE3;
    rom[221] = 120'h0DD300000000000000000000000;
    rom[222] = 120'h0DE300000000000000000000001;
    rom[223] = 120'h0DF14079D800000000000E00E13;
    rom[224] = 120'h0E0300000000000000000000000;
    rom[225] = 120'h0E1300000000000000000000000;
    rom[226] = 120'h0E2300000000000000000000000;
    rom[227] = 120'h0E3A43EB1909D00000000E40E93;
    rom[228] = 120'h0E4A43EAD091100000000E50E83;
    rom[229] = 120'h0E5041D8EC33900000000E60E73;
    rom[230] = 120'h0E6300000000000000000000001;
    rom[231] = 120'h0E7300000000000000000000000;
    rom[232] = 120'h0E8300000000000000000000000;
    rom[233] = 120'h0E9300000000000000000000001;
    rom[234] = 120'h0EA1408F6C00000000000EB0F43;
    rom[235] = 120'h0EBA43E00119700000000EC0F33;
    rom[236] = 120'h0EC041D8EC33900000000ED0F23;
    rom[237] = 120'h0ED1408F6400000000000EE0EF3;
    rom[238] = 120'h0EE300000000000000000000001;
    rom[239] = 120'h0EFA43DFB028A00000000F00F13;
    rom[240] = 120'h0F0300000000000000000000001;
    rom[241] = 120'h0F1300000000000000000000000;
    rom[242] = 120'h0F2300000000000000000000000;
    rom[243] = 120'h0F3300000000000000000000001;
    rom[244] = 120'h0F4300000000000000000000001;
    // Initialize remaining locations with zeros
    for (integer i = 245; i < ROM_DEPTH; i = i + 1) begin
        rom[i] = {NODE_WIDTH{1'b0}};
    end
end

always @(posedge clk) begin
    node_data <= rom[rom_addr];
end

endmodule 
